PK   �^Wڮo�  �
    cirkitFile.json�߮��u��.5�&���n�_��8 �I� �>�\�n��w��rK��M2V��Rif$:�ʌ&3������O����ؾ���������C����{���o�_���?���?�����i��������������Zڗ��-�{;�G_u�T]�tմ�mվ涞��m��������o�T����Grs�"������h3�_�߾�˟�������>M��m}5��Uu����e��?u{lÒڏf��������o���T����O������?�����u��?:��S����_?5i݇�j�9U�04���*���u���C���]���w]�|<w)�wd�b�N1��98� ��Sݧ0zO!9Oarݐ�1���u����+8�Nv���<}o=J�� ��/�����r|GǮ��$%`�⟲$����Y�~^�̢��Bd���"��?1�������,|ϭ�[�&�:M�:�c�W�s,yd��}�559�n|����5�'�'��$|wY}�I4ޓ�'�s��w(��9��*�<�O�����.N^����,���(N����>ͫ��"�L~^��t�n^����/Z�!2����Y��}n���o�����!2�	tCd����,����Y�k�"���N7D���k�"���N7Dfᯝn���_;����v�!2�tCd����,����Y�k�"���N7D���k�"���N7Dfᯝn���_;����v�!2�tCd����,����Y�k�"���N7D�1�k�"���N7DfᯝwcیKZSՎ}Wu�<Tː�j�z�e[��}矄p��'r��R��E���9������6�K��[��VuS	��U�����]۴�g���n����v���֮E��^Ms���ڷxA.;L�3�y�g08/�@^��'�x:�p��l���f6 ��e+��@�P�ܧs�._� �=q��LIԇ�e3���њd4��S����Le���5��,��Ż�2���i�����-�wmm�Ix�h	}�ݵȩg�}�%o��SO��\[�d4�ym�e��z���u��jjЇ[��]�����E=	�l6��Ҡ����m��Y7į�cN��l�}�%?�}۔���p��yRY��Nw=O*���Ie�$��<��D�2~����Ở'���篝n�_ۦ<��;�q3h/�U���N��.�U��7į-c.�^����߰����'��I������ԓ�?���Է	���]�����лkVSY�zw�j*�}��0�!���T~�p׬�����f5���0�5��,���YMeᯝw�j�{L���>����o���n;�9|&��O=	�s��Z��7MO ��U�O���v��^Փ�?�����*�C��Pe���u�,���.C����л�2TY�����QQ��o�b�E�mTT�պ9x��mT9�<@�u7�ۥ.X�9�<����e��z-�����*oa��h^��=U�1�jZ��j���I���.�EnY�`/�����-�}��9�����[}��V?�|8Ի�B�͠>�.�Fų�5�|.�:��]��4B�s��,�O����*���QRe��5J�,��FI��fp�騲���U^��@���K�b�d������G���Wo��a�l��\4s�{����}�N�v��Z���������w�~~.Y:�ѿ�H�{_���y�]����?O�k�TY��	w��*�<��Se�'�5z�,��FO���WTeᅸ�U����Se��Xw��*`������& �9\n#H�.諗>=���kzǧS���X��"w�z�S�Ӭ��K��M�'�^w��ݣΓ�zn��&��!;%�f��&�7�;��]~�(H���w
NA�ꮉW=	��殉We���5�,�����d��k�UY���]���o�xU~3x�ī�������]=��9��fr��{WR��,�>V����R� 9��}"�����z{�S��캽Y��u���q�_.�]�Γ�r盂��h��۩���ٽ��\�n���2�G '�����_���7�}����?��k�VY�W�En��>o��������������}�Mؼ�[ы;-�9x��ߊ^�p��q�"��y���}�"/���/�M���e�����T���������{�zwF����3�"|	l��p��X۽.�9�
 ϧ��Z�s��<]<����m�������s\d����9.��?�n�Y�t�{��,��m����Q�Ɛ�,�U�.:T�����.��v�Γp3������0��Bn�閷�wj�n�!��]p%���7mw2��Z���Ժ��Z�6�y����a�k����w�?����лݟZd����O-.��z��S�,��a��S�,�1`I�_�o��Y�����"�a�ݟZdᯝ��S�,���vj���v��O-�������Ņc�ݟZdᯝ��S�,���vj��>x�௝��S�,���vj���v��O-�������E��y�?���_;o��_x�k����"�ݟZdᯝ��S�,���vj��6x믝��S�,���vj���v��O-�������E��y�?����_;o��Y�k���MG�_u�m��w�$���.����j�X�Pv�eW4�v��.��ꏖծe��������`\d�;V��Ue�Xvy���9]d応G(?��v`�C�%�]�1�ڍ�v(�Ĳ�?&V���e�Xv���j7�ڡ���l��'�_|����]�w�LvE_O�)�hcD;#�%�%������[����/��ΎkX?����������
�/���.wX?ذ�����χ��M�/���/`�`��g��D~��$��������\hk|n�t��y����ί`�7��a�%�����j�~7��v?�~X~	�w~7���_������}q�Ǚ��Q�O/�9=�\�yj`���K0��;/X?�<�����B�6O,��;�������/��ί��ؾ��������/,��;�Ą����/���/;��x�~�}a��_�������`~_�{!��`���;�8�����/���o�a�`���K0��+oX?������>��,����v<H�8�?X~	�wf������`~g���?X~	�w�0������`~g�������?:�t��`�%�ߙ����_���y#�~��`�%�ߙ����_���_�B#��`���;�iX�z�������o$��?X~g"��?X~	�wf������`~g
��?X~	�w�G���_�ӟ�������������,�3���,��;��`�`���K0�3'�����u�ߡ9���y�_��]�����~��qCU�s���ɶ��� �5�_z��=�c��c_��_жo���o?�?���O�8t[_Mi{U�먫y��*�O��۰�����|T���H�����*W�A�Fս��@��;v8?�7i�o���|��hgF\����ˀ�{L鹪Z=uS���p�e@����ɪ�Lv8B;���R)����d�#����/`�=���Yx�s{�q��ʣ���J�dՅ);��v�Q;8G-znzƥ�Pe�g\�'�.g�����sԢ�'d���QvzB�:����!�����s䲧gH�,�C�-�ϐ�Y���{+��!!� ��W,?CBf��ϐ���/��J�|a���3$d�!��n)y�{z���<D~�2���x�~�m��,���;'9�R=_�;���lrx��>j��@� ���I�T�6O,?C�f�������x�/����<D~�{����x�~��b��9��`���3l�!��������I�T�6O,?C�f������/�~� K�|a���3l�!�9(?C��z��}�,������Y�����a�6����:���x�~��`�6��`���3l�!�����g�,�C�����Y������!`� ��,?C�f�����!`� ��,?C�f��?X~���<D?����x�~��`�6��`���3l�!�����g�,�C�����Y������!`� ��,?C�f�'�?X~���<D?����x�~��`�6��`���3l�!�����g�,�C��S`�!X�!�����g�,�C�����Y������!`� ��,�wA�����!0� ��,�w!���?d~R�ܛ�Ŀ��U0��u�Ѽ2֞��R5�GW�������������L��32���,�R���/��hgF\|�޶������eY����3���%�G\���(���<a�#�C�����ɪKv8B;���(���,a�#�C��ъ�ɪKv8B;���(���a�#�C����ɪKv8B;��o(���a�#�C����X]�(�C&�(?C>�z��O��
�TP~�|�<D?�b����x�~��`��	��`���3��!��v��g�',�C�-��0X������!`� ��,?CB`�l?X~���<d��,?C�_��?X~���<D?��?��<D?���}x�~��`�2�
��`���3d��!�����g��+�C���ϐ�W������!�� ��,?CF_ҥ���!�� ��,?CF_��?X~���<D�/����W�2��I�==C�_"?l_X~�"�ʇǉ�����T�`���3$�!����gH,�C���ϐX������!!� �v?,?CB`��2�g��~J�\����͓৞/l�X~���<D?�<���x�~����!`� я�Nv?r�_�l_X~���<D?ؾ���x�~�}a���`���3�!�}��Y��f�tv?r�_�$l_X~��	=n�O��K9>P�v?,?C�a��~X~�x�<D?�����x�~��a�����/�a�#���/��9�aOϐ��� l���A�|a���3�#�!����gHG,�C������xH�	�~X~�����W�p�4��WS�^U�:�j^����S���6,�����kp�K(0@��X��s�_�s^�/��u�ߡqܐ�<ׯ�q�n�u�����R5뜪n�j}�M����m���d�V";��ݛHH��N���p�v(�79���UP�p�v(;=|Q<Yu��Gh����œUN�p�v(;=|Q<Yu��Gh����œUW<�p�v(;=|Q<Yu��Gh����œUW:�p�v(;=|Q<Yu��Gh������,l,�pCu:[��!|� я�������`���3�/�!��6��g_,�C����X������!|� ��,?C�b�l;X~���<D?�z���x�~��`���f����x�~��`�����W������`���3�/�!�����g_,�C�����X������!|� ��,?C�b��?X~���<D?����xH��?X~���<D?����x�~��`�����6+���x�~��`��KO���`���3��!�����g�?,�C����X������!�� ��,?C�a�����!�� ��,?C~a��?X~���<D?�����x�~��������`���3��!�����g�/,�C���ϐ_X������!�� ��,?C a� �?X~�9<D?���	�x�~��`���`���3$�!�����gH,�C��?7����W������!� ��,?C`��?X~��<D?����xH��?X~�" 9<D?���{˺��~��QwK�5MWM��V�kn�y�v�ߠ9����!'���iyyܾ��_�,�9���ն�[ե4Vkj�*u�6oM���Q�O�������wx�;|�>��|���a�v�q��/9G^r�t=��}M�k������ۮ��e��i��--�1�7w�t�������K�_k/~-�t�S��^:�������ï�zm�x��s������Αws�k�_���^��Ny�1.Sյ�PM�����ꗡ9걻��ï՗�_:�Z{��k�Ý�_�����w�t��]/~}�k��;����׎w����^;�z�������fثn9�\ᵧjn�5{�����殗�V_:�Z|��k�ï��w*}�K�_�����w�t��]��s����^;�9�n�z����5�k��J��a�j�RM�+MiX�׶�������K�_�/~��t�����N��z���~^�~鏦��ט�j���W7�{����u��������]:���K�__w����.~}ݥ�o�sr�8�4W�z.2�sSe?PW�8��k��q4w�x��7�)��7�)��7�)��7�)��7�x��7�x����~���~��O���u�e�r�j����4U����4����t�����u��ףN:�z�I�_�:���Q'~=�ïG�t���k��n���3���2hL�T�W�4�ztÞRs��B:�z�I�_�:���Q'~=�ïG�t�����u��ףN:�fcm���3�z{�U��>|9��j�4��6�{w�z�~���~���~���~���~�z�~�z�~�z�~�z�~=��׫]�u��&���y���[�-���:�}[�F�t���^ƾ�����#O����en��M��Mz���{"���_����5�11��Pu�1W�:��9+�����_�����4��Tu۸��1���*-��5��w�|砕�o�}o�!��j��U�a�����jZ����i���ܕ�o|\פiʂ�c��]}�q�JN��l�Ż;w��_���ކt^���v��u�ex�M�n�t{���׿>-�k]�sJ|d#�6S��Q[�f��im��uw���7墨<	ڵ�_����jI�P5�<�ݔ�y���*���m��>�}��9W��ut�46{�ZS�׵m��8���_�p䪰�q2��2��93��9��إv��܄t����7�<���T�s�(4۫�ۡ=�m_C�{�+�_���MM���D���R��5�)����u>���S^:��;�e��-��DuM���s��|B���qjn�8��J��S��C5��9�#��:��ױ�c��=ޮ]H������z��W�o��5U������K���]w����&��.���}�/�Ԝ�
��c��:���:���_�۹��,X;�O�Tg隔����ݖ~mӼ���t��3nX�|W�I���r1�|x?��:�Gʏ�\3n�q��7羵�y�K�M�<h�f��>_�y�����u��YI��T�z�ao�<�f������^�֧ux�������*��(��i��`9�%�_�.�k�2Ǵ5��n�K�ߜ��''{;Uǐg]�g(k�g�mJ[����U#���_��}��=��-��6�:?��La������j#~S�~\�sN���1ўӔvJի����6���]:�fv�+bJ똋U��QyF���i��d����������eor�:ΩQ�������^M6�}���;��o��G���ўe�떧FK���A�����;w��;n�7i6U��ɔ��C����O�mO�w�r��ׯW�ïW���Ճ��W��v��u���I�1�����zMC:�zMC:�zMC:�zMC�ޛ�y7|��=z����r�I�9�:�3�ǳ"�c�mX�g��[�o��߾^�ӎ�^�ӎw����9�s�7�q�x����O��Z�-?���7xF_�:}t�z��������gׯ�_O���?�;����������������Ysڛ��<�n~^z�����*���{��/��g�_?�tP���P���*Tn&���ՙ�ϰ��z3�P��MH����r�[׳hq����Y�8����,Z:�f-！�f����a7��j�s��͢��/g�b-���H?9��q���y�z��sI��/'���w����I�?���ˉ���>�/�������4Z�u�Mw7�����9�����o۷?}��?���2�����_?�S9P��>_B3� ����3� ��&�@�Ծ������?����i�'�O�z٦z�1�SK� �j��b4R���8�ni}�&������_>F3�(}��4�����9Kd�q��6V�V�)���sB� ��ӋB� ����B� ���3C� ��ӇC� �Os����;/�����_��>�n��:������x���_�N���8�R}�q��S�q�e>G�89a���*6o�:N!՟�2'��7�	B�?Wp NR����p���ϵ"�6o�:N!��Oc���x���)�s�d�6o�:N!���b��:�bu�B:���8au���8�tn��q��x��q
��������ҹ�$�	��V�)�s[D�V�;��SH��}'���X���m�0NX�:N!�ۡa��:�cu�B:���8au���8�tn/�q��x��q
��	���������q�����qil�qIk�ڱ�����Z��VS?�S�,۲���"	H�+=�-2����"�v��_{܌���"��������+2�)����"������+2)����"���"��'��h�4z~ު��}�Z"��͕m�n�@*'�r�@*'�v�@*'�z'�|}E*'��}E*'��}E*'��'��'��'��}E����t:	J*��	��V�)���+B8au���o��"�Vǅn �Vǅn �Vǅn �Vǅn Վcu\�R9au\�R9q+)X������|��z1UN��!� $��H���v�t����"�ӄq��8�$����X��TNX��TNX��TNܚ86����"�6��TNX��TN�|\�R9a�q�H��q�H}����>Q�
�?��N��W�r��x���)$��H��ǅn �Vǅn �Vǅn �Vǅn �Vǅn ��9Vǅn �6�����"5;�R���\Y����������A@��$2��j�Hd�Ｂ�wWp�����O��@sz��U����������Z{��b�����6��7�j�Ċ6�$�����-t����-t����-t����-t����-t�� $)�H�!�g_Q,��*�E�U������Yƅ%}���5�6Ήe�q���.��vB��ʉ��cu\�R9au\�R9au\�R9au\�R9au\�R9au\�R9AHR_��	B���T;��ǅn �6��TN�JJK��9�Y��QB_���9�Y���C���v�8au\�+R9M�2��W�rUڙ��=�@���5�	����W�r����r��ĹEql>.t�������r���B7��	���@*'l>�K7���1���X�:�K71��TNX��TNX�[�SG�
}E*��Z���TN5�����r����r����r��U�n ��9��"t����8�$�eǖ�}X�f�S�CS����R�]��}=h}E����H���A@�>h#�	#H�+A@J_����A�A@��}������4FP-��� �ZڽL,�����I�?G�n
I�M��ne�2�V����DNX�Vv/9a\ٽL�!�Jʐ�	B���!�Vǅ�!ub�;���DNXWv/9AHR_��	����e"'I�+R9	�����:N!i�����:��^&r�긲{��	����e��긲{��	[GQv/9q+)�R
VǕ��DN�|\ٽL��Ǖ��DNXWv/9au\ٽL��qe�2�VǕ���EL��+�����:��^&r�긲{�ȉ[�ű:��^&r�긲{��	����e"'��+�����:��^&r�긲{�������e"'��+�����:��^&r�긲{�ȉ{�ɽ��긲{��	����e"'��+�����:��^&r�긲{�������e"'��S�@�}E��o�O�O�����V��۟�������5 ������5�p�3n��)D��)�k�ф�ڄ��5�p�?�]�]�r���Եѵ�5�k
��Ac�7���_�¨��C�xBt���B��c��c��\S��c
�u
�5�k
�Z�!��!�FpM!\Ϟ�c���|�n�`c�ްED2]A�+�v���c�R��
a�b؞��1�Ƹ��)���3�m�a�b؞��1�Ƹ��)���C��1N,�m�a{~��m�a�b؞ߔ�h��ް%�C؞���h��Bئ��7>!�M̛�7liXR�_�����)����U��AoĂ^����&Ɨ51�,�m�a{~�m�/a�b؞���h���k�!l�;��1����e!lS����mc|Y����F4F�_�6Ű=�u��6Ɨ��M1l�ovc�b|Y�����8F�_�6Ű=����6Ɨ��M1l�o�c��V��e!l�o�c���e!lS����mcޗ��M1lό�mc|Y����J��6Ɨ��M1l�̇mc|Y���̮��6Ɨ��M1l��m�_�6Ű=�Db���e!lS�3%F�_�6Ű=�]b���e!lS�3�&F۠/ɂ>%��e]�/�b|Y������6Ɨ��M1l��mc|Y����p��6Ɨ��M1l�,�mc|Y�����
Ѷ��e!lS�3,F�_�6Ű=3�b���e!lS�3�-F�_�6Ű=3�b���e!lS�3;/F۠�����_����>Ɨ��M1l�,�mc|Y����d��6Ɨ��M1l�l�m�:�o<�m�a{fd~aK|_6����)���2n�_�6�c��ۯN�_�QBئwlo/��6��T�c�U�0�2�������fٖ��a�^��b\�e��
kGu5�`vTP���Wo�.Q㢇�5��9{UT���aGu��j�^0.v�QA]�r%�k�w٫0*�kWs����q�Î
���+1^#���W��\�٫���;*��1�ǎ
�j\ذ���Fp5g��3��eM3U��1�+��={� ��6�vE��g�����X�����XR���֞�Z Kj�֞���c¬i��16,��={� ��6Ɗ���g�����ر����XR�K�֞�Z Kjc�Bؾ�^�a�71�,��={� ��6Ɨ���g����ߍ�����2k��*B�/ak�^-�%���e!l�٫���1�,��={� ��6��={U!ƗY�LUb|Y[{�j,�m[{��*B�/����"�������X�3)��={U!ƗY�LUb|Y[{�j,�m�������XR۠v�_fM3-�%���e!l�٫���1�,��={� ��6Ɨ���g�����������XR�_�֞�Z Kj��B�ڳW`�/b|Y[{�j,�m�/ak�^-�%���e!l�٫���1�,��={� ��6Ɨ���g�����������XR�_�֞�Z Kj��B�ڳW`Imc|Y[{�j,�m�/ak�^-�%����e!l�٫���1�,��={� ��6Ɨ���g�����������XR�_�֞�Z Kj��ˬi����1�,��={� ��6Ɨ���g�����������XR�_��m�*K&+�������XR�_��m�*Kj�ˬl�i_ڥߪ����ֶZ�~��~����ڦ�>�e��~gGUr7%Ts����x��Q1���U;*6�٫vTP����UQょ�5��9{UT���aGu��j�^0.t�QA]#���WE��vTP����UQ���5��9{UT���aGu��j�^0.l�QA]#���W��qU� �tl�٫�A�+�uٮ����XR���֞�Z Kjc�B�ڳW`Imc,X[{�j,�m�ak�^-�%���b!l�٫���1v,��={� ��6ƒ���g�����ز����X��B�/ak�^-�%���e!l�٫���A��b|�5ʹ ��6Ɨ���g�����������XR�_�֞�Z Kj��B�ڳW`Imc|Y[{�j,�m�/ak�^-�%���e!l�٫�dgR�/ak�^-�%���e!l�٫���1�,��={� ���+[�m9��={� ��6Ɨ��}��J4�[�LUb|Y[{�j,�m�/ak�^-�%���e!l�٫���1�,��={� ��6Ɨ���g���_����g��"��2k��*B�/ak�^-�%���e!l�٫���1��B�ڳW`Im�>%��e�4�XR�_�֞�Z Kj��B�ڳW`Imc|Y[{�j,�m�/ak�^-�%��ʖX�ak�^-�%����e!l�f���4SU�_�֞�Z Kj��B�ڳW`Imc|Y[{�j,�m�/ak�^-�%�����e�4�Xp�6��={U!ƗY�LUb|Y[{�j,�m�/ak�^-�%��y_�֞�Z K&+����o�W	_�&͔x�Y�W`���7i���1�,��={u�����R5뜪n�j}�M����m���}�*��q}��
���o0;*�k�w٫��E;*�kWs����q�Î
��՜�**`\찣��Fp5g��
:쨠�\�٫��E;*�kWs����q�Î
��՜�**`\ܰ���Fp5g��
6쨠�\�٫�>�pY�L�9|��
ak�^-�%��]1�˚fZ Kjc�B�ڳW`Imc�W[{�j,�m�ak�^-�%���a!l�٫���1V,��={� ��6Ǝ���g�����X�����XR�[�֞�Z K�Y��e!l�٫���1�,��={� ��6�X�/�������������XR�_�֞�Z Kj��B�ڳW`Imc|Y[{�j,�m�/ak�^-�%���e!l�٫���1�,��={� ��L��e!l�٫���1�,��={� ��6Ɨ���g�����+��2k�i,�m�/a�6{��%���e!l�٫���1�,��={� ��6Ɨ���g�����������XR�_�֞�Z K~���B�ڳW`Imc|Y[{�j,�m�/ak�^-�%���e!l�٫���A����2k�i,�m�/ak�^-�%���e!l�٫���1�,��={� ��6Ɨ���g�����������X���_��m�*Kj��B�ڳW`Imc|Y[{�j,�m�/ak�^-�%���e!l�٫���A11�̚fZ Kj��B�ڳW`Imc|Y[{�j,�m�/ak�^-�%���e!l�٫�d�R�/a�6{��%���e��UU�_�fj�^-��d�}��?�q���eN�0�C�m�Vu)�՚ڵJݼ�[ӯ�8}�JBP�EP:�GPeDP&efF4x�ћ�ᛘ��G��xmu�u�Pus�U���2�s��e<����H(��IBy�L��U�P/���\��*#�<V	��H(�UFu��eF�s��`���\e4����˱ԩ��q���݇jzu�\��W��Q��s��P����x�$�ǫ$�<^$	��F�UFBy�2�c��P��6��ˌ��*��0����h0�#�x�u?nG�7�^uˑ�D�=Uss�٢m��UFBy�N��e�P����x�$�=V	��H(�UFBy�2ڨ�/3z���Ì��*��<���_�0�UJm6^�XW똖j�_iJ�ڽ���H(��IBy�L��U�P/���\��*#�<V�yY��?�j�_cF�j���W7�{�̫0^$���"�<�	�q�H(��EBy/��x�P���r�:�4W��-U��M�mV]�㴮��N���
��ʙ��p��<��)(��f
�󺯂�0��y�WAy�Ť~YҺ�ղu�b��TMs���[׏}�0�PǮ��8v%�Ǳ+�<�]	�q�J(�cWBy���ؕP�n��u;�}����c��:���Yף���}���8v%�Ǳ+�<�]	�q�J(�cWBy���ؕPǮ��F���~�i���{�C��R5G�yǽS�W��*�y�JAy^�RP������U�y}UAy^_UP��W�Ǳ[�^�2�s56��(�Z-K�f�>��u4��cWBy^�Xƾ�����#ς����en3JS/k�^�!��P����ښ�T��e��昫e��꜊�G�ʿQ?s�P���3u���q?�c��6UZڱk���YX�PP�u��qȃ���s�x��j�뺚�iyu}�ƵtQP��tפiʚ������)�=k��k�W�EBy�R7{�鼾G�u�P���U��ڛ�݆I�EBy�2-�k]��M�	��T-��R3�˴6��t�P���vy8�k��^)�t{��y��i��nJ�B����<���h��:�\����U����kM�^׶�i	�ː�#�-���y���4�qNk7v�];��I(�s�>�s�tTC7���y>�l��o��طu|I��((�\�nj�&?��,W�6��yN�^Hm��1̇p�$��{��u�wcw�:�5]�8s��|����qj�{ZAy~l��7�P��k��ȵ��C�u,����ʺ�����u�{=�ǫΕayMպ�Z��m��j���x�P�����j�哙�>���Wzj^�^x5���uJ�����ȥo�f����t>fS��mR~��v[��M���EBy~Nk�o�<�ٗ\���Q���֡>R~��R�<��g]�65�y����w�����+=��ju��SBy~�Ӹ{S�Y`v|���}���>��+���3@Ay�Fk��)���_���F��<����1m�k�#	�Y�#���v��!O��6O��.O�۔��u7��ڡ��ȥ���k�<�Y�|FC��;�Ώ�<!���8�]�u���h��u8'�[��j�97k�T�ک^m�Q��"�<ϥr�Nis��\��#O��<�O]�K���(������ò7�b��0��3J�Tӫ����u����<9�ml��<6�Ǻ��ᒲ�G~���n]$��{z�� ;��?��G~�x�	���O�'��'�VP.�kA��Z�����c#��Z���f�(�kA��Z���$�<�i������f]��q�|������y\��`W35f'f'f'f7�(n��kN}�)Y��(�ӫ�V̯�x|���s�IO3l��Q�˫�=0����]l>G��L١y`~��>zN�eFq�<��i�ܵ��v��#ۮ����f�c�$��K(��Y���<�QP�g5
��FAy~$((#rF���y �:h�2�W��H0ϳ	�yV#�<�j$f�	��¬F�z�(f5��(>�i���R��qW�J	�s/c?v.6��x���o<0��x�e�<0���8�ni=0��x��W{5q�`�_�����<u�Q��Y��������ǿ�����������Ӿ��o�O��e��a?���>̦�iY۪}�m=OC����/�~����?-�k�V�D��.a՟30�T��FP�93DA@��,a՟3V�T�~FP�9�FA@��aտ���Um�lcu;a��B�12'�v'�xSH�/����p
����1����"N!տ�R�V���SH�/����Ϳ�	8V���SH�/�'��7X���_V,NXo�:N!տ��0��:�`u�B�Y�a�8V�[��SH�n�'n%�[J��x��q
��������ҹ�4�	��-V�)�s�b�V�;��SH�.�'��wX���]Y1Nܚ8�(�����ҹ{&�	��V�)�s�F�V�;��SH��ث���X�����0NX�:N!���a������M���X���]�0NX�:N!��"a��:>`u�B:w��8au|�글4�͸�5U��wg��P-CZ����k�m�^R_�������A@J_���jϏL�����  ��Hd)}E"#H�+A@J_��R��DF��W��H�jse��B7��	��B7��	��B7��	��B7��	��B7��	��B7��	��B7��	��B7��	��B7�:�����r������B7��	��B7��	��B7��	��B7��	��B7��	��B7��	��B7��	��B7�jǱ:.t���:.t����n)��B7��	��B7��	��B7��	��B7��	��B7��	��B7��	��B7�����q�H��q�H��q�H�ĭ�s��X��TNX��TNX��TNX��TNX��TNX���W?X��TNX��TNX��TNX��TN��M��&Vǅn �Vǅn �Vǅn �Vǅn �Vǅn ��9Vǅn �Vǩn ��h���]����ܿlm�e뇪��yi��m�N�+����"�ѳ�"#H�+aW���)2����"�����  ��Hd)}E"#H�+A@J_�������Um�lcu[�R9a�[�R9a�[�R9a�[�R9a�[�R9a\�R9a5\�R9aU\�R9au\�R'�X��TN�����cu\�R9au\�R9au\�R9au\�R9au\�R9au\�R9au\�R9au\�R�8Vǅn �Vǅn ����-�`u\�R9au\�R9au\�R9au\�R9au\�R9au\�R9au\�R1�:.t���:.t���:.t���5qnQ��B7��	��B7��	��B7��	��B7��	��B7��	��B7�����B7��	��B7��	��B7��	��B7�ʉ{�ɽ�����r����r����r����r�����0����r��8�$�-S��}X�f�S�CS����R�]��}=h}E����H���A@�>h#�	#H�McI��i�  i4�$탦1���}�4F������AK$W�����me�2�V����DNX�Vv/9a�[ٽL��oe�2�V����DNXWv/9aU\ٽL��qe�2qb��qe�2�7��&�XWv/9au\ٽL��qe�2�VǕ��DNXWv/9au\ٽL��qe�2�VǕ��D;��qe�2�VǕ��DN�J
����qe�2�VǕ��DNXWv/9au\ٽL��qe�2�VǕ��DNXWv/1�:��^&r�긲{��	����e"'nM�[�긲{��	����e"'��+�����:��^&r�긲{��	����e���+�����:��^&r�긲{��	����e"'��&�z����e"'��+�����:��^&r�긲{��	����e�s��+�����:Nu]���ۿ�?U?-���7[���oZ~������� ��fPS�µθ��]#����G�k�k�µ�hCtmCt���B�f��k�k��5σBt�Ct���B��9J��C��\S��c�u�5�k
�ZL!�N!�FpM!\�9D�9D��)���cbW����m��6�uٮߕb�W�q^!lS۳�<F���6Ű={�c��q`!lS۳�?F��6Ű=�a��6Ɖ��M1l�o1b��qc!lS��mcY����6&F�W�6Ű=��y���Bئ��J1�����)����U��AoĂ^����&Ɨ51�,�m�a{~�m�/a�b؞���h��Bئ��7�1�����)���me��1�,�m�a{~#�m�/a�b؞ߺ�h��Bئ��7�1�I1�,�m�a{~{�m�/a�b؞�P�h��Bئ���1�u+�+���6Ɨ�1�,�m�a{~��m�/a�b؞1�����)�확�m�/a�b؞�1�����)��]�m�/a�b؞!�v1�,�m�a{f��h��Bئ�g&J��1�,�m�a{f��h��Bئ�gFM��A_�}J�˺_�����)���m�/a�b؞�G1�����)����m�/a�b؞YT1�����)�황�m��Bئ�g6X��1�,�m�a{f��h��Bئ�gV[��1�,�m�a{f��h��Bئ�gv^��A)A11����e}�/a�b؞Y�1�����)����m�/a�b؞ْ1�����)�홑����Bئ�g�g��1�,�m�a{f��h��B�&3۱m�%��jǾ��a�eHk5�S=uͲ-��Ü�jGŸ��W���̎
��՜�**`��쨠�\�٫��;*�kWs����q�Î
��՜�**`\谣��Fp5g��
9쨠�\�٫��;*�kWs����qqÎ
��՜�**`\ذ���Fp5g��3��eM3U��1�+��={� ��6�v��.k�i,�m��
ak�^-�%���_!l�٫���1,��={� ��6Ɔ���g�����X�����XR�;�֞�Z Kjc�B�ڳW`ImclY[{�j,�f!Ɨ���g�����������XR۠Wb1�̚fZ Kj��B�ڳW`Imc|Y[{�j,�m�/ak�^-�%���e!l�٫���1�,��={� ��6Ɨ���g�����������X�3)Ɨ���g�����������XR�_�֞�Z KjԮ�ˬi����1�,��={� ��6Ɨ���g�����������XR�_�֞�Z Kj��B�ڳW`Imc|Y[{�j,�eC�/ak�^-�%���e!l�٫���1�,��={� ��6Ɨ���g����}J�ˬi����1�,��={� ��6Ɨ���g�����������XR�_�֞�Z Kj��B�ڳW`�/�c|Y[{�j,�m�/ak�^-�%���e!l�٫���1�,��={� ��6Ɨ���g�����|��2k�i,�m�/ak�^-�%���e!l�٫���1�,��={� ��6Ɨ���g����J1�,��={� ��6Ɨ���g������2+�mڗv鷪?��ꦵ�������黶i�s���j�^����o0;*�kWs�����沣��Fp5g��
<쨠�\�٫���;*�kWs����q�Î
��՜�**`\䰣��Fp5g��
8쨠�\�٫���;*�kWs����qaÎ
��՜����c�5�T���X�����XR� �㻬i����1�+��={� ��6�~���g�����X�����XR��֞�Z Kjc�B�ڳW`Imc�X[{�j,�m�%ak�^-�%���e!l�٫�䛅_�֞�Z Kj��B�ڳW`Im�^���2k�i,�m�/ak�^-�%���e!l�٫���1�,��={� ��6Ɨ���g�����������XR�_�֞�Z Kj��B�ڳW`�Τ_�֞�Z Kj��B�ڳW`Imc|Y[{�j,�mP�b�/kc|Y��B�ڳWUb|�5�T!Ɨ���g�����������XR�_�֞�Z Kj��B�ڳW`Imc|Y[{�j,�eC�/ak�^-�%���e!l�٫���1�,��={� ��6Ɨ���g����}J�ˬi����1�,��={� ��6Ɨ���g�����������XR�_�֞�Z Kj��B�ڳW`�/�c|Y[{�j,�m�/ak�^-�%���e!l�٫���1�,��={� ��6Ɨ���g�����|��2k�i,�m�/ak�^-�%���e!l�٫���1�,��={� ��6Ɨ���g����J1�,��={� ��6Ɨ���g������2+�ejҺKլs��ah��56U귣붽����U;*�՜�jGu5�`vTP����UQ��eGu��j�^0.x�QA]#���WE��vTP����UQ�B��5��9{UT���aGu��j�^0.p�QA]#���WE��vTP����UQ��5��9{U���.k��:���\!l�٫���A�+�wY�L`Imc�W[{�j,�m��
ak�^-�%���`!l�٫���16,��={� ��6Ɗ���g�����ر����XR�K�֞�Z Kjc�B�ڳW`�71�,��={� ��6Ɨ���g�������e�4�XR�_�֞�Z Kj��B�ڳW`Imc|Y[{�j,�m�/ak�^-�%���e!l�٫���1�,��={� ��6Ɨ���g����I1�,��={� ��6Ɨ���g�����������XR۠v�_fM3-�%���e!l�٫���1�,��={� ��6Ɨ���g�����������XR�_�֞�Z Kj��B�ڳW`�/b|Y[{�j,�m�/ak�^-�%���e!l�٫���1�,��={� ��6�S�_fM3-�%���e!l�٫���1�,��={� ��6Ɨ���g�����������XR�_�֞�Z K~��B�ڳW`Imc|Y[{�j,�m�/ak�^-�%���e!l�٫���1�,��={� ��6(�#ƗY�L`Imc|Y[{�j,�m�/ak�^-�%���e!l�٫���1�,��={� �LV��e!l�٫���1�,��={� ��6ƗIl�o���o?�?����i�v���ߪ.��ZS�V���yk����AIJ���J���ʀ��ʄ��̨�/3z3|3~3���^�5����n�nn�j���Z�}���>W	��:I(��IBy�J��E�P�k�Xe$��*#�<V	��h����}�23~����8��z9�:�U;.Sյ�PM�����ꗡ9�{�2��u�P/���x�$�ǋ$�0���H(�UFBy�2�c��F4x���\e4f�>W�q������fثn9�赧jn�5[������H(��IBy�L��U�P/���\��*#�<V	��H(�UFu��eF�s��`���\e4���5�k��J���k�j�RM�+MiX�׶<W	��:I(��IBy�J��E�P�k�Xe$��*3/K��GSm�k�(�Q��<V���zo�yƋ��8^$���"�<�	�q�H(��EBy/��:^.QG��_���ֹ��ͪ�~���5��8a�WAy^9SP����u3�y�LAy^�UP��}f�<��*(����/KZ��Z�.W̶��iNS��a���OCf���ؕPǮ��8v%�Ǳ+�<�]	�q�J(�cWBy����m��n��ϓ���AqL�T�W�4�ztÞR#�o�PǮ��8v%�Ǳ+�<�]	�q�J(�cWBy���ؕP�רֶۏ<5��W]u�}��c[��HC?o�w�����B��</P)(��S
���򼾪�<��*(��
������8v�׫]�u��&�e^�e���ҧt��f�a�J(���ط[_Ws{�YPߴմ�mFi�emҫ=����#��]_[��jS�U�s��s]�S��h^�7�g.��:C~�u=U�6���܆�JK;vM=��8k
ʳ.{;y�U�v.�\�}]W�:-��OӸ��.
ʳ��4MY�}�P�w�8e��am�u��
�H(�\�f��!�������u]�j^{Ӷ�0)�H(�\��~��|��#;ᵙ�%�Uj�y�֦�^�.��{�.��v���+e�n��4U3���Mi��Q�pPP��u�X�VǜT�:�j��z�)����6�=-�<r�p�b��a6��;�9�F5�i��.�k'x5	�y���{n��j�\��9χ��U�������!	����MM��Z�������9�)���ua>������|O���n�\'���gnR���w�:N�rO+(�πm����q|͹b�v�y轎e���QY��P����q��<�xչ2,��Z��T뗵��\͗^/��5�\��|2��'�7�JO�+���X��NIY�UP����lsִ���l���Mʏ���nK��iޞ�H(���am���>���Ԕ2J?��:�G�O�\��紂��֦�5/�4�8����|��u��C�n�A�cJ(�πz�ao�<̎������^�֧ux����]x((��h��>�v�K>�5׈u��\@��8��y-�}$�<�r���N�1�	P��i���It�Җ���]Y;�P��Ӿu힧=��h��|��1�'D[�G��NBy~M���$u��S�=�f픪W;5ëm2�P_$��T.�)�c��}�KU}�	����s�~�垖P�{zX�&W����zF�jz5S��|��5�P��/G���ў���X�<;\R�������ޭ����|OϹdgW�����O/?a�<���������

��q-HBy\�Pׂ$�ǵ 	�q-HBy\�Pׂ$�ǵ m�A����]03~��`4f'f'f'f'f7�(n�̌��3�f7�(n�Q�0��aFqˌ��yO�8�k5��t�G�]�>���rlÒ��y	���|C)(�����|;)(�w���|3)(�����|+)(�w�4��ˌ^aV#�0�W��H0�f53��Y�ÌbaV#�@5��¬F�aF�0��`�Q,�j$f��ˌ���j��?������}�ӷ�>����?�������O��~��O˶�>���Ƿ�^�O?���׿���Ӿ��o�O��mڗv�<��n���������黶iϤ���I���cیKZSՎ}w���eHk5�S=uͲ-��·��r�����������[��ｿ�� �8�`r���$�1p��!�b�����J����w9�.6��� ��d&���%�j�M�^:�J�K��k���!/V�XMC�i.k�H��ͣ�~:��=�ӷ>:���zչ��O�vp3������K�����97iݳ��97i;���A4�>��A��N�+H���݃�ղ��{P��aY���U���ӽ����e\���@"�\�7�!1�婻v��n��D��ʓ�Ϧ��Uq��i�
7H#��n�b�_�fu���|<J�#�N���ҽ�$�:I���{;�G_���4]5-�}�m=OC������{6��(�t5��㵑#�5Nq����T��e��}��}�(f'p��Uד2���m���
\�f�����t5'	\����^� ���x9!_��*����*,�y�����4��Uep�|�2�6�*���&4pݢ���*�M���_�Xv��Dh�*��Nu}u/��;���g뇏�uE��W�@�������>����*�x|ׅ�2p�ěz�2p�񹬉*���nގ��si��~�2�ߍ�z����}=������LUD�r��	8	�ށOF�C�����t��'����}����R�*�[�3����v?���!�O��yȾV�=������~�wk�i�]hu1K7��ד��u�����M��_���$�Tn�n�ߌq����������}�>��_Ǣ8�7������2�h�oMN�����K����ޞ@N�����R����98�����}���ɗ'���s���!o�v�➧}�j���ѥJs��@�e����+m��[߯_���~}���eC�����J�����7�R�����/��?����s�]��������)ק.fe9~;ON��~0���/��Ǟ5��������Y����������������������������_�����`)��?_
�ᏙBhiS t
!BdO1D��7D~�$*�H�p�s�Nx<ÊN�bX�aU+<��aEGWݗ��+�
a�Y}��;�׹�ߙP���o�-�"Ɛ��4��"D��?�R����W"�I���"@BC*c� ye �������%8�Z�#b��>.��:���v/��0[�!D���BK9�n��a��q](E������"�� A�}@6�
��CX�I}�Vt`��-����!���>���ǰ���~�wـ*H� ��Dx 	�� B�Dx�c���{���"��,B��� ��!2D��B�W�[ ��Q/��gE�����?��a^%C���$����]��[^��ύ ڔ!$�2D��S��w�bO"D�)CA�4He�� � #!Bܻo=����Q1��XF�Ĩ�#@����|䢧�o?��|a��%��F���]�U�񖙉��� �; 8�[�A?
y#<�<o��!ҽ"@��"oY���"������E ���w��P�����
�P����u<�2��Q�O����uAp9?�,�/�g�Q޼)-H3���n���ހ�7$~ߜu?!8n����gD��Se8�ݯ���'�$��� 	>;@�iX i�  �`d��9�w��;�=s�!+����㷏�y�y�����;�_�?~����������Q�����l7D��~n�|�Y�!��~�����Io;�s���8]��_r|��������Jo;�p����+)ץ8ݔ����������]��7���	6��������O����I�d�����G��>'&~n�̣x�1>cq�<��٘~n��t^?7Ƨ��21p���sZ����N����A^�a�����G��˨,�%P�?1����%����7_�rN���S���@O� /����/,]���e�'���p�7���z*K�	����C�� ���pc|�l�y�1>���<����~���
��!���q���ۏ�	��̸[���1>��<�z��ԏ�ٯ������~����~����~����~����~����~����~����~����~��n?���@=�c|�?�y ����>C��<�z��ԏ�����PO{���12���12���1�>~�PO���1�?�PO���b�;-�I�~��gq'�����[��>y'���bk�+w�;y�/�\;)����$�uպ�n	�'��/�vm��n�e�Mn��r�q��������e���S�����������S� �T�뗈�M�m�n�v��<��}�i�� ��m������M�vn�vۼ�o���nr>ao{Y������܉E�p��ZΧl���Ɠڵ�د�,�)�J��P��t�Ԯ���}��A���C��F��q?Ư�(^@o�E7=%*�R����<��|��� j�m?��(��� �W��m?��(��� *bE��~�_{J~���������K��q��Cѹ���2Le	�b?Ư�(ߩ�\�z������D�C�-��yE����u=(ܷ�'*�p�6��<��}�x�� V�����yE�L�oOT@�m<Qy ����0�m<Qy ����D}�����e�������\s�_[[�c�\y��=4����Zܿ��:��A���bTZofͮթ�.�P�o;\T@��pQy ����E����u1P�o;\T�D�����%�&�y!�d� J?7�}�������ݓLdᆨo�XDn���kEd�x��һ��E�\vBɁ�_8����%�\� �y�_8�v�x��r��#��~���*�]��eߍZ-����x�Qy u���E�T���P�o;\T@��miQy ����E���x�tQy�1�6����6��!J�H�����|��rو���a�z��t�l ң���t=��F�\6ި,�	8P�o;\T@��pQy u���E�����P�o;\T@��pQy�1�dTn��.�:����0/��pQy+o�����ef���#m����x7�{���h����T��M3�w�N�p����I/޼k��nh�/����neؽ�Xt��7���'��G�<!n[iTĪ7��̸o[iT�����F�̸o[iT�����F�̸�7k#�U�7�����7k#�u�7���'*�7}7�E![+�����zw��t�}7*�7sy�ܛ��ڡ�;He�u��]�{��㜝�_���.�
y�=���~���������Qy k2�=;��r`M�gG�̸�=;}?Ү��DiG�!v��X�!v��X W�6�Mcᆸ��Y�!��~Dn��������,��t��F���W�7;z\��k� ^�k�q��z�H�!��\oR%V�7���Z�,���f��='DZ@��c<m�$� ����K"�\�o�$� 
���K"�d�o�$�pc��q4*7F}�?�� ��m��:���ozg�w�i��t>0���|T��tMf�uTZ@-~���q�v���]�D�@�~���s�q��H(���!�<��}���(���!�<��}��h���}���X���I�A�Y�@��I�L���Cy ����D@=��I������D@=��I�������e>����$� ���~H"����$� V��e`����$� ���~H"����$� ���~H"����$� ���~H�����$� ���~H"����$� ���~H"��b����!�<�zz�������!�<�zz�������!��^�zz��������w]#��o�O�O�����T��۟���������q�g/^��%�_�Y���/���֯��c�%�_������~_�}��c��9;X����`~y�q���G��B��C���8����̯�a�FX?�_��������K0��c���a�X~	�w�V���/���P��L8�!�U w,�e�=mZ�Zm[`��fxv����f�h�g�0�!�W`��fxv:��&f�h�g�6�!mT`��fxv���ff�h�gw<�!mX�2�n=l��Ii�h3L4��#��U���g�i3<�����.f�h��� �������b��4���&�����!�b`��fx~Dk��#|��rNT`��a���ihS3L4���+ZC������r�֐650�D3<�z�5�]�0��/��Vڶ����ڐ֐�-0�D3<���5�m�0�ϯ<i�1ڶ��/Tii�3L4���ZZC���0��/�ii�3L4��fZCڧ����"�֐�)0�D3<�&�5�}
�0��/�a;ڧ������֐�)0�D3<hi�3L4�3=�֐�)0�D3<�h�Z�Zh���>��}
�0���ZCڧ���L�5�}
�0�ϤZCڧ���Li�5�}
�0�τXÞ�)0�D3<�qhi�3L4�3ه֐�)0�D3<S�hi�3L4�3Q�֐�)0�D3<Ӡh�/��O�i���>��}
�0��.ZCڧ���L�5�}
�0���3Z�/.�m�c�T��-���\��	��8|&�$�p�	��u�h�3Lo�����/��1�q�oo�ީ���ٜ�����f\Қ�v컪�Z��VS?�S�,۲�>)�v<�ߛ������^vxDN�~��!r��ބ~wy�R��ӗ��x��,?C�x��҂я�g�W^V��!�}���ۯ�z���9�;"'��:(����`�C�����x59��#r�v<DN��!�P<_y�������葮��S^`��!r�����\��2z:[~p3�j�� ���3�����IX �hH���%�� �ѐ�20CK$a �!��I��2�`��?��i3�D 2>���p���������S���ВPX �h��gZ���v4z��zʴ���K(�5�'Ss�ʮ ���65z��zʴ��Z
 ��&�C��%�� ����80CK`a �!�q`����@FC���-	����,CKB�zʴ�����S�M�ВPX �h�2�$��L�=�O=e���-	��L'
�ВP��2m[��?��i�3�$ 2��b`����@FC����)z�_ �!�S`����@FCڧ�-	�����O�Z
 i�3�$ 2�>fhI(, d4�}
�ВPX �t|�>fhI(, d4�}
�ВPX �hH���%�� �ѐ�)0CKBa �!�S`����@FCڧ�-	�����O�Z
 i�3�$ 2�>fhI(, d4�}
�ВPX �|JI���%�� �ѐ�)0CKBa �!�S`����@FCڧ�-	�����O�Z
 ���i���� 2�>fhI(, d4�}
�ВPX �hH���%�� �ѐ�)0�w�  YB���%e� �ѐ�)0�w��  �!�St�۴/��oU[�Mk[-[?T]?�K�wm�vo��=�x�Q��m0��Ǎ|y��[���x ?C��ϔ#(��|s��9Y~�A�|� ;��ϐ#(��l��x�~,?Cp�x����!�������ʦߎ����3$��+~;��ϐ(��l��x�~,?C4�x��ѷ�!���р��Wv��̄�eh�TO�$�)�]	�ВX �hH[��%� �ѐ�#0CK` �!mI`��,�@FCږ�-Y�����5�Z��
 i{3��� 2�fhI�+ d4�m
�В�W ȬT�>fh��+ d4�}
���W �h��2�}���W �hH���%ϯ �ѐ�)0CK�_ �!�S`��<�@FCڧ�-y~����O�Z��
 i�3��� 2�>fh��+ d:Bh�3��� 2�>fh��+ d4�}
�В�W �h���o�go(L��W �HJ���x��^��j[�|FR���-i������Z��
 i3��� 2�.fhI�+ d4�]�В�W ��3�����%�� ���65z��zʴ��Z��
 iS3��� 2�/_`���@FC������z����m�Z��
 i�3��� 2Ҷfh	�+ d4�m���W �h���ws���3�F�.FO�Ofh�TO��)��,р����Z� i3�D 2�.fh�, d4�]��X �h��O�=x� ��b��(Lؒ�*@�=�O=e���-I�������Z� �w10CKR` �QB��Ụ��2Ԝ)Z_c��K���Ц&��X���=*p�߻�A��%tp�����R5뜪n�j}�M����m�3��7����M� ���'�Qv<D?�ߛA���Kv<D?��!8P<_yy������3��+/���X~��@�|�e;���(���`�C�c������я�g�W��v<D?��!8P<_�����X~��@u�K=�O���fh	, d4�m�C�X�@FCڊ�-�������Z� iK3� 2Ҷfh	, d4��	��X �hH���%8� �ѐ�(0CKp` �!mS`����@f���)0CKp` �!�S`����@FC��	�S�X�@FCڧ�-������O�Z� i�3� 2�>fh	, d4�}
��X �hH���%8� �ѐ�)0CKp` �B���%8� �ѐ�)0CKp` �!�S`����@FC����)z_ �!�S`��A@FCڧ�-р����O�Z� i�3�D 2�>fh�, d4�}
��X �t^�>fh�, d4�}
�ВX �hH���%� �ѐ�)0CK` �!�)
�S���@FCڧ�-Y�����O�Z�  i�3�d 2�>fh�, d4�}
���W �|�H����?�ѐ�)0CK�_ �!�S`����@FCڧ�-i����O�Z��
 ���i���� 2�>fh��+ d4�}
���W �hH���%ޯ �ѐ�)0CK�_ �$B���x?�ѐ�)�~�Sڶ�xBb���!�}��?�q���eN�0�C�m�Vu)�՚ڵJݼ�[ӯ�8}������y|�<�s�;��Ǐ��'��w���w&�L�1���0݌�u_�����ơ�涫�y٫e��~K�x��]������7�@:��
H��\ �x��7U@:��
H��T���*��� ���*�x��]� nF�V/�R��j�e��v��սrA�^�24G=vwU@:��H��\���+ s����T���* S��o��6~��;婢��wU@���k��q;����[�<�x��c��ck������7�@:��H��\��� ����
H��T���* S�����xW4 �����(��5�X��fK��u��i�����4��k[t��5������7W@:��H�{�����7U`^���i�[w+ɍ4_��b�)�_��=;�5��c��!��-l�T+���5���e���y�IUf2I}I2�^�
����fd�c0"x�����t�񋡲��J�N�sf�h�C�����#��G�⏴?�i�?��,/�����d#�J4�U.� �Ԧi:K�0�h^�ee�XR��d�XJ���X^��m�X^�xT�5mZ]խp��SKME�j�Ԓ*�B!�� �� �� �� �� �� �� �� ��x�n��&;ތ�ie�*ƚf���E�E �� �� �� �� �� �� �� �� �X.����FڎT�sa|=�u���m��E<���2!,���� ,���rq,���rq,��G�G��׺��fT:~�Tu-O:t��:�?�?��Z�V��������Ԗ;~F�ю�)�?���7]���ax�*�[Ս%�踐�u�v{?��݈�1�hu?��ܗ���5ׂ-�����}ϵr��l;���U#	�Lc�NHjt#�ߏ���?��1Nk�v�� #~�q�4�am�8F�⏽�������6TBpU5M#�Zu=�U&�����&]���\��0S��e�֦a�t���c�a�yJ�7U�u�񋾪�U3���Pkk�F�c���d�}S֙��2��U�PW3i΢�⏼_Q583�:���~:Y't�-m��7"@���W�^b�P)�����$X�U�+>�m�;E��?�y��q����8�ɝ%��:$S�z������c�o�uӻ�#g�Γ��V^�F������L�J��:�58KF���n4s��x�⏽�tO��;��oݙ�i��!놓���ZF���_3g'�ݎ3ʒ��3�sH��PKI(������%���Nk܌�%N��A��x[ˆS������?�p�E�����~����U��@��H|�C�c��r�:[�^�~�*#]��F�n� �QQ���_bt�zV9?��/��n�]�Jڨ��6}��"�1�7��ơf����q=���v���`Z��Q�C������sSʹ�;'�Ν䔶N������y?1}+x���u�+�~�Ĝ+��~d�?���5�n�t�=nh�q�TǙ���?�83Ii�����28ױw�,Ϋ�Ʋx�����O�=s�k�'�:~YW�c.���k���!���?�V���\N�u�SM�7�6c+���C���g]�uqJ%��4�RW����\�l{���#��?������rݶf�I�:�Q]$;�G�$;�G���ᙋ���e��S��9�EhX�VA.Hi.Ji.Li.NY.NY��q*mN}>N�ɩ�7�R���[Z��/���S9��i������>�S���#9�pn�`�V��m��spAP���1u�C�j�$C���y2̓A�7<�Q݆'���b���w'��Hu��زњ�=�T���/��@���\�F��\�FȨ��4��@l�4Ǯm86&4�C��vׄz�>���@��;6&4�C�mX␣	��;6:�hB����9�а��.��/�W_o����W���7��B�~^}����l#Fx����hbG�=~⨶�)�p��#)i�H�L��W�&���Cv�|�l���E�/��U����*B�m�
�a�З���YX��Bd�̮
��/_*Q�UY0 �K�j����d�ŒX �`@V4,�%d�����_0 ��d}�V`�{	`�z� �,/E�������d������t�R$`�q�`�p����-�L�-;0��V닓^�� �R-�
d�J����td�#9ة�l�`#9���F6r𑃟�|�_���	�|�=������q��@\�?���m��k���u����I��G�����gmͤ���G-���L;W�:WP�qHr#�����JV�u�ݐ����C3E2y"��X�H*O$�!�I�$7D!��:��~��7�P2W���P�� �r�
u;P(gW|�t�P�f
E7�2�fG�ABћ�A�Y���L�TA��/%���mtOJ3壤��t�[P�+a�&�[m�s%,��[F��L	Y�V�2~T�J�JJ�6$�3�k"��3߂^ޘ1޻�)Ԇ�FM�k
u׶���Bez�|�cc�޿ �Bm�,���"G(������|[T�-M?*G�\ن��� �T�<��-�CT(�)����*�d[SA�
������rͻ̌��F��rͻ̲�tSS<׼�PD�
��)���1�4Zb#:�y���FŽ_�_S�K���!�.�_��5#��y���������4��y� Yu�җ$	u�s���8�˘�L�^�;ˉ5�s+O9�mQ�����h����/�08T�o`�*d�%	����L�#kOBD�7�s���[9@�B�0*�Ƹ&��(S(�/���Sp� e
Ŝ�L� @�h�Qeڈ�Ep( e
�� ��Ԕg��M��E�Ғ9n�HP��ֵ!_p� E��+ې0����تl#Ɠ����BtT��hX�x
�A+���\ϲ��vZX�x�e)�欝�6�Y��T��gY#�������p����H����ɜ 7Y;7���#c^4�2�b���i$��?k���`���\��*˹w��EyS �0!���F���ͩ�x!���������h��[f�����(8K��rρ�O��+��͝��)���/eQ��vug��􅤔
Fz(�I�_���Ү��H�������%�ǚ'�K���dh&�׿��78��*2����|q������z֋���2'p^��k;A!�]_��Z�H�9밾Nؗ.8%��U'�}؃/����0�m���d	L�cmĤ�f	����p��(8E�	���%P0'N�mI����Ym��Mм��+��h�&˦�Ѡ�6��	�q���SV|qT�89�U8�ٞ����O7�b?�[�����7W�~3��z)�~�1��_��_$.E�/��"��K����H�E�Rd�"{)�^��A}u�gu����>��:)����F��:���:��N��:)��Z��V��:���za�^��6��za�8���&�0_/l����&�0_/l����&�0_/l����&�0_/|����'�p_/|���;��>��z�^��>��z�^��>��z�^��1�E�z�^��1�E�z�^���lY|��I/�׋��"|��I/�׋��"|��I/�׋��"}��I/�׋��"}��I/�׋��"}��g���EN� 7�a�v���t&}��I��׵���|��I/�׋���|��I/�׋���|��I/�׋z�6�a�v���t�|��I��׵���}��I/�׋���}��I/�׋���}��I/�׋���}���A�׋���}��I/�׋��b|��I/�׋��b|��I/�׋��b|��I/�׋���������Ǜ��{{7��|�}|�D��U�q������Fs}#5�`g���~xrB@i�/uUL�A˲2��ڠ4â�UM�NuCY��W3����1��,������O�q%�<���������?���ӧ��cP����p{7f���������?�O��Ә����~�|w����������t����o���c�
����>�6���������﮾yrҺ��S}�y�ۧ��CL�9�a����~������Ə, ��������S�w��k�܆�)s����i[�*#SI��R�U�0�$}7�S<q����r�����í������	`����҂�q�>�R)����q��E6�%H��u�`s�0�
Kx�.&g_r~���IZ&?��2�I�U��\2̥\?���>���sw{������b���ܸ���v���2����~�l��>�����^𩉃IE/н<���TE9��aļ�� ����:�q�?{�LD�x��F����E���-�-%�����:��ԅ�s�6t�)Է�ε�z�^�l�T`gݟ��e�l^��%r^�f%��_�G�f�l;��Iҭ"��a.�R���U�w)A���s{t�/Ի��t G�N�M��TD�\<�%�\�N��hۉ>m;�c��]+���wm�0s�0�
s�0׶��I�s��I�?I�5��7q�^ܺ.g�[�tŴvA9�]�XSW�m\���'�l�K�H�5.?��9i�����J�E_���+#C�ì�ͲP�R�5F�˹f��K�k��#����"ȵ=�m�誗�;�ڊ��U�������"�a#�AO]F2���*���E�k���-Ug$�ɭ<�� ��,+C��^Wn.�Q:r������Z=�D^S��z<��5��ϟ�.RlY=_P��d��d��	|%a�r���o�QrrKwn7�ɣ9�Om�I6�D���ư6�˗�N�dk|̅]��Ĕ����Ś���w,	���e�1�K��(		�z b��s��.�8�r"�8e�b�\Om�Y�X��LŁf���*�/ B�$�`>W��?ޞl��v��G����=;���g'������;z�k���y��G}���prmǙ1k�tHs=���`�r��XK�����"��/>���H�F=�N���N?��������l���H�ȩox�^����?5��o�4��w�]��oM;�r!��v��޿���������f�W�����q��sIjY��B�ִ���MX�lK˙E9y��WMe>ˍ`�H��􃖌1N8�����
{v�'�^���U!V^�)wQ,ג��j�ra
]P�T.�|7�_!L���q��B%5�J+�S�Z$�|aM��5��`*H9�����$����;4�&hr�tM����Q��,7ss:=�c��¬.gN��Ah�9��R��g�����?|�^xZF���{��;�9DY5�b���kM�f��ҟt��	�����ݿ�*`�v�b��Q@WH"�9��ɡp��������"��0@w�Bӫv��s����C t�+� 5G�|G@Y�� ��!����P�� �Ve��p���P�� �l���s0���r6@� �*v����9X-|U�u)�mm�E?8H�n�\������պ�����Z�W���cFV���r��EtE�i�h�ز�Is�V%jZ��.A^p�{��L�<�Ë�q�I�J��VB}e�����n4s�ip)'�s�/�L�{f���̤��2�.�=��wDW��Lմ�T�n8�����ǡ@fR.���=i��A��锑�N�kfk#����S�\����:6����߉�	̋P���1���������"��ֺܲ���f��Q�9���;�ֲ�Զ���H%ɗ����py�ZV��j�ye������R�Qd�F�����E�*��~�����ele�����U��P����H�Z�F����7
\�~����A�5��rxM����{ճ��W��֢�ZI�сۦ�P9I�g�뼇;_.Ŵ~�.�U�M5�^U��.�T����Na��=�ky��x_��⒗�����ཨ�u���E<DTF��~d��-�q9_�.ޗ�}���HWf�z#io��Y;\6�:n�+%j=�e]&.'���z��_.�\�O��ƨ6R7j�@�J���q07��a����N0�9I����Nޡl}��;~���c��ԍ����$��%Ce�����qm���H���_;~���E�+[���J�{�H�_YW�c���uV���$�~/E���j�{9��8~ہ��|D���M�WuM�1X:4c�A�;I��ߩ�~�%�[g��ՒrH��k���U-�\���PY�\�:aHϙm�C�.�Q/Gϝ�R.�:z.��)H�E2�5U�d�z&��3����ߞ^6^U��˽~��}���/ ��ȟЮ�N��9(
)�\�%���mUָn��/Zjq�{g��A���1!��t��-�ȼL�y�Ћ2�(�2�x"s�����I/��L��Q���	�Ο��L-�Ģ�/�袌�˄��	�(;��t>tz��22/�|���erQ&��޻e��-Y�^	������gx3ú��c��T"�L�Yr�Y��yS����r���aޝռ������`f� �%r^��%fV"	�>�RB�d|V��y�����P�{��w^5�חϾ<h��GW������O�K�.��:�|�o�*=������������o���Hj͗��f�Ǣz��n��=����C�����?���'����;�������o���/�]r�����u�����ۻ�w���{B�kyȍ=���u�ڠky襶���?�(`�����ﰠ7d���^���jT�q������ӷ�ӏ�������_�&�i�v,���4>��~����y|~v�n�_�0R\o�Y%Wd?����/"��ܺhs��[��&����+��!�32���<�(x�q��ǁG%��tl���Y��Pa0�_xdQ����#��N�<�<h�ԯgآe�C�����C���dd�b��do���=�ѥ�>4��=%K  Q@�t(J�� *(1r ��Iк� B��!�"{S 1Z@�8 1z �h*�$ �d3���hri�O�?��C}��ͩ����������������_D���]te-�Ӓl<��͚_m~�Jͯ�7���# 5���M��m~�J�o�7��軛_b�/=�OI���� @Iyl	�� �A��@_k��[��B9���B��(@_k��[�� � @~=`e�Z;` �~w �!����,�kA� ��wC@`I�?�(
z��&��a��������?<u��.3�Jn7���R����/Tt�G�d{���Qs7Pv�4�(�(K�h�K�!��E�TA���L0�7D)n����N�����u�R�k2A?0�A������@e���������|�:K���5Y &��m��X�q�\�{�a��s�T1>
2,:��m����G�Q��$Q����j!_jE�T
��⬬������q&˘� �4G���"��e��c�g	�����"<��!�n���vP��avI�55�gj䁦F�4SC9bB�M�
J��t4�e�&��؁^����`FMU<,��M��V�0�|���N&:�ڎH�w#�o�ؼXB��!������z	486�H�Z��F,�������e⌚Er@PlN���d�}��v��ɥ=ΗIL �,J�K��$�D�Ƞ�����5�U�2��c��@x%n�������<?d�lҸwH�G�v��Ϙ�J�a˧{��߉����D`��������d2�V�i���/���vT�^�TF��پ���x��f�oM�1p$���� �^T[��ug��i��VP��"��2 �)��9�4�!ˊQ���̄�D_	/��e���;CXS����YDԕ`LT�v_�;ˉ5�s+_8Sg�B����߃�~��;�c�Ϳ� ��bW���/*��-�wB@`~�Gv�+~6+k�|%�����{�A�
xd����g��������@��2E!+����[Cj�ѦWu�K+���N���v��%Q�c�b؋���aI��i�ƕ=%��p\Q����i�?���[*e[,�q K�U$�E�@�%�0������ �����Xʎ"X҄�\T�",0���
��'P�)t�-�`�l%B=8��֍ 	h�H[@rp�]�`ДE ���!�&�X1�`f������9)�QA��W)
h�57�7��
 �C�Gx��C�U�2���D=^�k"W' A�hnE�����
P��~!��W���������w� Z>��׏���dpu����N$�~' �K�⯷�@ 2�0p��ä��aQ�_R�V�vS͑fE:t�J;����{�ЦJَ�z ��#*l,E\�U<Юg�����ུKَ�z\���#��X |_S`͠�Nf8<����OG0��~m-��l
�_Mp�_�6�a�y�E�܉��H��y��[����xFe-O�=T���yF��P)��!����;�m�as���8�9q2be-B!���$�JQz�Gl�G�7���m��#�2�l�f<����/t��p:oٯB��O��������
��s�����V�D�ݹ��41��C��I�52�nCfu�L��6�0*��c��Ҏ�Mah�<����Jz�u2��i��<h����CV���iMZ�W��������S�:�"�	Y��=�0]��h�FZ'Bt����*y>��X<]��?��j�$�;I��hЊ��`��!����{���)��5BVg���ZZ�5h���U[Z%o�&i࣒h�l�u���1�c��@��� ���S2�0z
�&Y0A���-��6���ߚ���^���U��r�v*#,�q�I�D봺�<h��t4p~��bad��������~
�'[2!���;��BvguI"Nڧ������C�:_)�]a�S��b�5]��xYq�
�N�������COa�d� &hu8�=��V�`��G{Of��sZ6�K:��@�)u�nݘA��m�q�0�=�6��v����8~
�']2!�#�=��Q��5h��Pw��k���`�R����h�H�}Z7f�>����ˋCT�uz} ���)G���)l�T��ü�5]��P0/����;m�1�j�v�R']o�A^�v�U�N0�u��;��z���~��W�'�o��U
�N:+"zA8�uV�e`'�Ѱ&+x��~�R���Rpب�(��/���w�a��w�����ƕp@M�xت��xq,"���;^����� C�o� ק'y�	��D����� ([.��k�c�T�)FUi����$$򍄋0n�Ɏ7���q�ت�D��!�U�nH���&�k��ZUJ��v��X#C��f"?ڠ��#����
F�;>�#�{{��$j��4
D�buJ���z�n{c^�WYP�.��uX[�.���W�2�}�8$�z�R�V�Fh� ��
�/�gь�J��2��*���u�+��k��U5�ECǜ}�P��/(�H!�#��
�`�c,�(e����>S��z�m�И葅������hof�b;�2m�-�.=&n��hښl@�< H�کa �v�<5�[�E4H'-AF��1K�Cֽ��b������d��g�����Ѝ[�wޱ6W��ܽ-�tK(fiT%���ag.\B�Z�������@T�5/�*pI�RI��b�FU�z?�m�Z�&�[M㑡t(S��0�b��ޖJ��4���i�u00BB՚,l�G����d�Q=yuoS%~��YWI{O�+��jM ��vNxd �j-�(}�%��j��YQ9K�*鼅u� #��5����p�iC�a�"���/�t�3*gi�$�0g\a���,da��њu�{c_�;%�������Q9K�*�м�s�0�՚,�!\��@\5]����ӝ����B����*M�R%h�}�f�<����R�>�ܠi�)�򦱳��6��v'M�bI35�� D�Y���. ����ۏ�4��~�n돏Wߌ�y<=����C}�������~����8~��\��� PK   �^Wġ�e� M� /   images/ff07c967-2774-423d-b98a-e9b309260373.png�US��gpwwww��K��������=��a ��ð�V����[_�K?�����Qj_�P���   ����  ��o ��'3�� ��m�����)Ԝ,m~Y  �9i�j�:��W>'�P���=
���Y(yxbJDE��Sis'�Jp4S4[4C;��r4C��e��H�3Ӂ���@�����ϻ|~��i�M��Mn2 �*�BD�<ҥd(6���Ig�$�e �%䳚D��d���~���vU7ڟ����h	�< IZ@=qjF�Y���v��օٵ���@�r"�&�����(�X8l��]����_�<B v���_y�F��V� ��z���Xe���/����M��߀��ߑ�h�=�ٱ��p-�潔>g����IlٺC0��86�Eߓ��&P�������`C�s��c�L�����aE��#�����94�GL���˵A��#�#�
h>�^�'n6�H>щU��X��#Eǂ�9�x�"Cꫥ��_ RN�3����+�6#�����\jۮ)N!K�j*����uz�]��7�մ
����8��#�$�R_gP5sL��~E�̓]��ء��}���X��F&\��}�5�0�L}N�7����60��;�́������
(tQ���Չ0�
(��k�,��BLk�p�\���s"�I���&q���I=��1`�$i"����%�(4w#Ƃڨ������j����;HY��d�P+�*��"0γ��&�d�R�!���f�#�����$v�HR�Ҧ�p���j��/�N�
Rf���a�"�%�Q�	e�Ahg�t����k�$��)�,�l�+C������3C+;]�$��	��Pӂ{u-���/#��j���+I����h)RkSw^�8�&�)+̴fn� ;,n�e�;�M;�>�s~������7s���c�(���☌s���A1�.����D��A}Ъ�/&wBwRw�VL������G��ih��]g�/����M�z���r"�umco{{7���^� � � d�@rZ5�Q~)I	m�U�U9k�M�{l�(&�"x�d���J5;9&8Y�:�نMAf��{b|"[��B��Jsd��|�:�+�|j0}_����mDc��\�����o�F�L��Z��y�4�K����,�ٿMk��+���T,�R�F�F��� T$�٠�����N���A�����ʨ��J�5��S�%1�hK����f�f��f�t{ţy͓�������Y�Yź��X-L-?��Mw��	�	��bgN�N�z7x���>�q�t���y���r�~�,����ي-K��XO-�V�(�-Ϣ��<��r�O{���YGز/lW��������+j28
�Nd�^����sI�%)��W�'���Ӄ��K��9]m����� �`��s/� ���Z���B�JF��������wkI��_��m��aIXN��}�16��eָ\���Qθ�3Ӽ}�D829�2Q=z/��c�gٻ�^�k�<�T��i�յG��<+*�DHS���P��w�i�r�r%˄���x������m���)~=���V�o��H�۫z�wU�Wj$�Z����ͮ8B���NE�S�g���Kk#:��;"Ǧ��;�Cd1�Hf5f�#��΢���X�.~o]j]�\�o��p���8h�G�Ϙ%Dl��d�tlh^�^��U�x���^�>�g7i�E�����+��s�`8�U������W����������|�}D@�@��� ����#u�-��v�m�Rd�J^��D��S�Q�'.�]��e[�g��ȉ��:K�G��q�N ����ۯnVv�^fDx��R�}!��$?�5I�Ie�d���w5��  �	��UΣWm�t����=�}]}�����y�=�xd�����"ײ,�z���t��@�D�����N���?l"����úJE��0
�@�`�0�"��O�^�Y�Z�%P�8w�ؿx��nSh�0:o6O�}M�HH?R���ɧ��0y�-��D�j�yb=��5}�Rz�Q��X������Mr9�,S/�������ҷ��}��͞'y�3����g�F=��>#yi���ivU(?pkOg����g��=8���Z�^-W۰.2N���Q�D�R�R����\�V�|2�64�z�ܴaI�]�ؘ��g?{>���?i�����,{�;n��R�{�=�թ������l�(5�誉i5d�`�ۖݤ۠�C��^�o��{dOcL��$�bؾ1)7>�1��"�t�T��»�\î/�-)�eww�ܶz+zr{�|�ժjm~<��	���pcss�oA��qf�qH�����}(OV���Q�}��ϕUl�=֭z��憔ޚ^1���Teh�q�6�=�6E�~CwKO����D��kU�c�g����Zw��Q�4}�������y���ˆ0;�Q�����04���	�U�.�[���w�G�*+����S'mعӹ*���͛�=k�Ug��uzGo۽�>G�[�]�ŝ>�S}�W��"}���!����w�&di"eblE%�w`��ۅ�ޞ�|Y�ձ+��Gr�W�|��4�c�EѶ ���ׇ1^�F���h��G�?,��?>VvWw!+�+f�=K�]��{]�I�I�W��	�/�_n����g8��e��*�BZ������̰�R��
����kKq@� ��H1�}^N������l<�ð<�ASp��9 *1�$�	wo����Т9�޾ޟ��h�'<�t�
��K��<_�B����I�� f��g�:O   � #������oݯ��CDVf'E��6ϧ/�<�h�D��ߐ�$yl$C�0Yu����y�%֠
Q0e0�'~lVi^�+����:~]�}t�=�=�֝��F�I\֟eE�Ņ`����������?�?Ї�BݭKy���竩��ʐ�*J��8����̧�X�[��0�t�XW���L��/N�����!S��#����M�|"X����̐��ϫϵ ?�UH[���˹c��U���G6�̪i��y�ZR�(g����`�T���z��QĮ'�Z��zJ�C��C�U|�J|	'�uuM9��9�T[[���9�5avwFP�s��;`�ͅ��cl3"�J05�:=�/Td�x��>5[Cb���n����v9��ב_[��a?�q�3G�e�h*������K�h�������d�3#�;{h���u7�ŀ���+U�����)�<>�e:3亿�<�EǼ��uէot��k(�!w-_W�|R�f���5��[K�V��C�7��Dr���2��	'���w�y�OG�σgn.�+tu����Cv�^�ZcLj�kɅ�RLjuN�{�Oz櫘��
����u�#F,�"/w�iO�
�?�����s�m|N|��tCN�7�?�DL���MȆy��zew�ކ~���hpp�PgJۣb2����v7C�vv�4 �żt�0�3UH�G���,Q^�	
^�&�(t@⧬m�^�.3B�C���:�����|DU��j��:z�<:�$Cn���*<,�P��݁ݰHd�Okg�9f�O-�j�^ �b,&+���Ó��>�ԚY?��G�u��Q�m�C*�Z��"2��8�/�2��lK�q�BmJ[����SK�In�i<��:/T+iM0�����VG1/�;)��dH`\� �[�c��2�<�Mp�<Λ�� �����n�&�������'�-<zbb�&6�@��u`���Y7K_7�>x[n�%c�6�VR^K���e"�l4�U�Y[Ӏ��
�m]dw��s[��q�Ξ�9c�� �{s��q�&�c{w0��qy�a���y�2���H��w��]�Ŭ��Gv\DGl�u D�՜G�>����M����b���x>Y��=���ث�vM�ZId��	aQ�ii}�a��ӝ��"��(���b�AT��Z>Jhװn�
��q� �t�3
��Vӻ����P��G�(E���s����t��{�K&���������];aV(�����Ox�v��0��=�]�)�Na_��ծ$,lg=��D�K���}�Q6Q�Kv�]�n[T�}���&[G+�>78d���`P�%��rOr皀���n������sߚtU)�T�@՜�6F5&7��[#dH�u�N�i81Kzc�O�E4_D��ڴв�ʳ�?ovn����,�-��][ ~�M2�s��N� spz�t~�ڽ]�4�����7��a�C� ����}ҡom:������ǃ�ˇ����ѧ�މ]�_ߺ�y�T�+��Kx.��e7�N���\����nA��+�
�������Hdv^�҇v���eYU ��O�p�~����u�R�,�s�\T�������d��_�XN����FD��%�;	Zc�p"�_J�C���5A�c"���͡Z'�N$:[5$�,*�JA �� k���5�+R{���&+t�	��{�g�M*aRۨi�}k���9���	j&�.M�����0�~_Nc���,�I;�K�s�唞a!E�D��Cf�Mr��8nLu���41��� ���� ����b4v����]��e@6>�٤���m�8�������^p]3]���G7�������~K����4?��?�6���{0���ʗmҁi�[0��z��2c4�,y!$G;����L(��:�0����se�D_[o��EN\|e�Y3�j��ᓤ,�6^h�_����\ne��N���Ǻ�3{OM@���`~Q��Zĸ�ɺ��3����0)�r5^n�7�r�Ⱥ�;�|���+�*�7�extuF龍��L�
�n5J8^���|��3�ϒ3�|sۯ�Pwn���_��l�,�HR~`����?�::�%�։:kO�c�
c��j�Q���GV4�˺\V���@7��Phihwc&N�/?^��~��_��W|2�ɂ��.�E��s�S^^���Mج���=�
��n�蝳�M��qF����$����H�����q1\$W��oZ��w98<�[��A/jc�h�5=�+�ՅC�1/Y���@i����x�E�oS	K�@B�|��:!�@�Sg8M����^�=��X�*�ԩ�4���l=���ʚ�Wqq"0�DB x]�w3t(Vڳ1i�$���\c�;�Q�+���� v~$Kac�������	s7�(	 ��@��� ��E���{_�s;��EcG����@Ǻ�1��z]Kp+`��O�Z�zR.3vo=�h���d/<S�Fo�ӽdg[�I�<���iFn���S_&P9���W+z	��E��P$B'��]�>��~�-�Y��D&��R�񸻴�0� s=+�P����K��A���{Wz�E�ˍs\�Fr`�O|`о��Iѷ����i�\�?��?�`����*�Y����p��<K��� }�EM���2�wi4A�������o^���F��Z�/nw����5 �L'���M�$��\�C��f�%^"g��X;�����Hw�4.��e�x!������5�X�x-ئ�("S��/vB5�������1���G��ؐ���~U拰X'�L��\i/��#)�#�RB�ю������{Mm�Ա{rZ����l��N�m.���B_Ö�gu���
'I�:�)^���������|oI&��=H�x�L,��J��?w��x����=�:��vF�c�u��l���$c�������4���N�`�!���Vp@o�L{��1)l�.2���9��z����4��me�����$k�1�ت�9�sxxu��ql���^�M`γ h��d9M��6 �9�Il��U���vx:�u�������
v� =�s���H�T6�#�C���n?"�|o3�l�j*��h !�OX�t����]��G|uV�L�:������(��`U�8�{F}@��3RP��0q�]l,�X�РιV�r^�I_���U$!���� �W��)��7�ˮ@�3�	��a��A�'���; q�/<h?ev�U�`mme�W�u�w���a*�H����w�h��R�H���z�I]��s�9��uR.y�V�DNӲ����S�����/L(td�[0I�/�Uo!n��i
�a�-x��u�S��2(N���̽�i�=
v3�6۠8^�x��.���W5/�:�њ��&bsU�m͑��|PH�sn�B? j��0�ӭi�u?x�m��-�\�|�&�����Sf�Q�,)�:��kT<�o#�L52���x��n�U	��QI�Re/$���Q��64�t��l<��ǇRf܄ϯp�
���8�W�T�WݡU���~�qӾ^��$�f���tb`Pu�"�Hh�9Li1y�?��0�
Fm�w$���J~%�&Vy$Sd�l-K���6�:G^�;����Cc��m6�.��o6|T�x��յ0N-;����A��xB�T�x�l8��J�Ku�In����ޘ�Q�)y��2��]hն&Pm��x�<��9
����"7��"� ��|m&E`[�ɞ)� qCc��|E���{�,���^låz"B�V��\ 0���fs�ϰ`�W��<�{"�ǀH�����9��p�gyw��237_c1�I�=����;ۣ́@S�)°ȢREgtB��2�O�A�W,e�gz@���rA�~�����˜հ�UVC�_���op�/Gf�7#��YhA���هۀ��ܷ��0�*�T^����n>��ΧG�cH�(��cc�1��8f��5�E����,s�ɯ��-�!Ƅ�Ą1hϳ\��˜&��C�Fo��c�;�
#�*��;�i���[>�ߟ[��&�G��Ȫ$&���Hm;�x��h D�I�u�'�q���YZ�Vzv]�NkQ(%�r����WI
(�3[)��ف�?�):��7�#�1Ƥ�*�D���N��#��~�Vn�`]6�/�䈽�<�����X�7��A���uћ�J��fH��[M(�G���vD���^��4c�0�c�a�;�36*����P���-J{_I7�L�Fv;bv����kF��y�=G�Ջ���|�hq��娃�������t�E�d����=k>x'<�R�
��
��_��=�-�.����������:i2��p�u�,0H��+�>I���D�qpm�Q޲ۆv?w�|��M��<H)b�B�r�9!(���F�k����C)8~�C[S��=˥��S>vn<(�����S��܇�����OF_&�P�~|*!�_��#�z�.�^r���cx�Z)� X)i�Қ"G5��4Ƭ^X��.g��~1i	h���2rV
����L��?w�f�6�\���I���m��s)*m'�X�+,Z}�(�������ؐI1��N�o�c�����y�b&�P���K:#(�i(���؞��w�t������������A�o�wI۾�D�.��]6r؈�H<��6��<�>�_n�,��<�\��w~�C����U���p���X �@�D�������@u��+�*܎{,�{��L�G�ó]��*r� _&��@HE�=�NJ~M�!�l��&JD ����{&�8v�'2%�~�K>Θ(�ˡ��Oh��@Χ�L�OK������t��lF�|��bip�] �^��3]F���W
�v����-9��'�˶�ߥߍHGV1Y�C��9��x/}�>|���}	��h2�Q��1#�  ڮ"�>j5���y,�mS @Co5žC�kP�M�����G��Oe�Y�ޖ��7�ڊ�5�;'`J'Z�46h �����:Ak��fgjOT�MN���Y�/�����|�hr�$g&�ۃ��)��L�����bJ,��tN]���Z��
���v[��Z2�'�!	��c�DLH{�{Ϝ�� b�R⪡�������OPM�q�u�RKD�qzl״�����n6S�Ƶۗ�|�="b-M��%��k�g	�A2IE[�6���	)(�r�>'�#z�Q~h���ۘ�56Pb��"� 3*�L��~[�h t[�^f�~K����r�F���D�b���� /�3�p�	�aP���ii�<S<��p��� W�ڲ��$:�ě��i����<D���6AFX��)_ ����z	h_w�[�3o5�~�?/�i�P˩	����A}���n��@T����0��N��?T�}����P�bx�\����3Q�[����q�]/����O+�}:�¶$�a��z �U�Aߗ�`���1���Q��B��j�{���̵��K;=A��>�7�"l~[��ZUfR���6���B	���-�q�ZvIww�N�.ۤf"X�����Bf�"p<�3%�jO���`�U�2v�	zm���hǧ�_�#j�|�6/x�%�Ro�8؇w��}gY�3T����d���碶�(.���z���+��7ӷ���M]l�c>�DJrL؎p�1�
�0���O
�J�Hb�zȀr�z�2������-m��t}��_ :��
���u4̹������{���G'�1�zϡ�ؕ	+�F��p,�>�!A����-\4C���xأ��������OPqr�Dp������>#.�'o���5�%w����\W�j���/4��N��b�
��;����7��w�-Y�O�b��|���gGjS��-6yt�ј-r�/�� �Ym��O��~�����N�k�Ï�l�/1��k
���ۼ8R������D�T�=�H��IZ�w\��]!����s�%��I_��qA%�|��~��ƥ�	��o�	M�.)Z�u�BM��X|q�e���2���l��i��^s���څ8R8��i���¡�5-���Vȷ��{�jOt;P��y�>x:s�2(���&���@h,�Q�{������b��<�[�we!i,��&0�J�B�N@E�ld�������S�Z7��Da�6��9���BY�~6zU
��,���XI�0��,&�`w��V?��K��9��-���٭ :�"�rP.��v��N���7�k,��&2��g�b�m�h��궃��~��k��\�)ǌU8�T��Hx��є��,�~UC���	Hň�:��UN�3�@�ʔ)4c��9'�����]��B��<g� �*(�h�0�S��x�B�
�]�T�(��?:])�L�����H��.�2�.+$���p��"`inu���5����@��0�aQ�$�̪m_���zH[��dS<hɺ���o��6Ղ�@Ҍ�I�B/�s�eX"bߖ��j�7+$�~�kٕ����vG}\�/|�<;��͘���m4֪������a�r��'F��.T�hcoy�����E��� �1_���	��V��YƐiy�H��c��&�:�<�@�� -\jYƔ������a
6``"��R{�X��t��"��"�D%�A���{. E�k��O�OP������ �Wa��y� Ñ1��*]~���.l����w��@������92!{ZG�-��
�6�]��=����T�h��";|��n�'���2����t|���T�v[e�8x��U��P����o�z��ѩ��Q��F0h���]{����������d���ZW���^�w�~�&B�ef��?t���-�,Y��kQ�-w��]G���r>B����5]�����h�ͧN��#����o���"�b��,t�:�����1�;�O-=v_Dڑ��h���M�ߌs��)s���dڸb�+6i8���K���jᝡ��Lѹٗl��R��N���,�p�<���jmDv�u_pݵs�U��jz{PgԭV�u�a���K��A��_w�S���뿊�������I8J���1��HD���'�R�����گk��`܊���� ���R��<Ago�k����<�F
Կ�(�2LV��̝��J��s��,�f�X���M���� 8�L�V2�)�����{ي����)D(yn��Ȯ!�5Zc�Ԣ�x\{�
��&#(��5[T�n��<���zD��<Z�	��1�E#����J�z��ǒ�-+������I���>a�X!�y���I���&�l�>m�ۧ�G�;���Yvs�:�!&P"�b�G\֢G��[uS���A�{�EX�T
�}� "5�y��������K�?�a�M�l��j����6;@�V�6���8 ��/O���|xm�m)���K.�M�!� �#��򫼹6���oN_������i o����!��OO&���緊��ė#��u�w+B�w&/���^���^���T��O�w%��m�~�K�pBݐ ��UZ$`%4���<����g.�����؆>X���we�H������ZK� n��;2�!�I/h
�V~�E콝&��f�c<�o�V���[ �:e$��q�0޶�&�/�!L�!_�2��<�쾙�����'I�j��~C��1Wp�F����+�㚂�S�66$�}]���V��]<�S��m����G��E��&K�I�O��\SZ����3�r�b��:Ƭ���_�2Q\D�oCx��\L�F`�ЅR>j_1����v�����4���e=��<���`N���L�[J1�*����v!�xU��F�l�'������ȑ� �t�%J=�4I����b!��[M�R����YS`4�S�c�H~u��7�bs1��ȿ
� ^��g��
�=�cf8C�3�a0�noGҶ	��������PF~	u���>��nE�t��`4YcZƕ�-��~���1y�ڤo,�P% F��<0B���g;D����D�Eݰ����QO��:�{'/�\`����c�LhQ����dq�\�<9�����R[[1�If�Lb��y�`u˦��^��:/ݨů���^�ڣ:���E�@�&p}5����
.��Wel�tf��A�bWض�-W��o���!�d���;bA�ܐMc���@E������g�����W�X%��2+Y?E/!�׏�Rt#��~�}��kȈ��z/Ll|}x�gYѹL*���3��3�|��,��/ܶo/�{��F�����٢���%� �x��zE�p��73-�և(zAvz�-v�1e-^�O����C��O��#����c�m�@'j�.���tC���v�����Ynhr��/J��t/���V�sm�1j���g�?�7�Q�'D��4�0��:H	�_���C����%���,L�g��7��n�0�PU
��Wq��:��rG�����*l�����tČ�� {T�G��24D�ţ�7���;b�Lsꕒn�|z�~>�E(����76�K������#Ra�w@� fn$,cҏ�Uqa��Zv�Q�s\�_'aҐ��Ū=��ɤ���8�%�C�J;��������4�A�{'vm�ӳ�Q�1�C�/���A�],S������=�i=�;)
MC����[۪����=2V
�׽�&kX�b��b�/�zx�΃Yk�XJ1��A�6ѱ�3�A���m��F��A��eve��2L}׭\��V#?���L����	/�,�i��:/�4DǛ#�C��>�{WTƅ�ǣ�!�d~�{���C�&��`>��Ϻ_|�|c̸��?x���؞��V��4d�y�mh
����y�f�WӉƔ���hkDer�Y����f&o�ڟ�e��ù"�8�����Y��-Cg�-4������<��*Ŗ
Bh<��0fy�r���*`�lܺ�Lݵ���EYR��������=DBż�1f�����b0C� �ռ ��\�K�@D��,�;,�>G�>_�'{J ��"o���<�f�o+1�W	Jk��mJdw}�<\_^A�=���h�W�U��e��Vpy?B��,���.l�<�9N���n0c�פ�Eup�	�=#��8�4�2T��3L�zV*C펵`G��8�s8Q���N��^0C#��#��nׁh��[r��"?,fL9�]�;�=���h�\���������9�aoQ����#��We��~�m�o����;J�7i5���֮��#�����"��A�<�|�_���XƓ�>V�]��n,y6H��8������l�d-m7��S���ԅ#���W�v���;y��|�2��yir�჏�c]������|0K����5M:�o@"�ܙv�M��j�h%,���]�����~^�?�$� ���n�JtaW3����v�S�����W�&�T)�<c-�U �k��XJ&����=>q�j`����Wǳ�=`�	U�sW����a�4Ͷ�c���|��g�k����J5�qèV �Z^?N���ܰ����u*��e�<9���o
��䫶Iq���o >vM/R�1���8L���2Z�8�w��fr�xn�nb����>�	+C�g��	�.N���Sb���pi��?��y�d��-1�ڣ_��D�7�R��K���yM(�SEdiAE_�f�~ߺ�X�S``��-p��XE��#�±`լ� �S�`��M��	�"��C��/��dXޚ�!�{c2Mh��M�)l]���><;��Fk�N�� ���J?|�kJ���B\��f��i/yV� ɵĖ�q��g�0΁\������Nܮ�wA�=�����!8偡�aq��f� �j�6��<�H�6��>�U�Аq��5F	QyVr�V�ߒ�Յr7�f,lݷ�:�Q<���hW�ߩ�~6zm� ����i��0�Ė;)��~V�6'l�=��X�ᶉY*7����QmsD�u¯g���@N��ɖ�o���b�T�u�
ߌ�/�����d�Y���/�3Br.�^�,.dk�z���9Ȳe�;��E�&���%�-p���������8}����_eůD�Z�_F���)��'Iה�z��##������
R�	$";�b�^l��XL�ۄY��+ų!\�9U��ꪥ�"�x]���q�zzP���0r�I���c/�.�(a.��f��6���K�`P��t�$��j)+�$�t�����q�#Cc�a�AT\��x��`Y;"��!�V��)1�E�<gNX�J�\?{�c����/��s"$�MwP�zH��e�z���u�}���rk
Q�vs��}���؂"����<�ҽ6������� �꣢"q@<J�5������H�$B���iǌ[�pF�L��H�s�g��l�Ccߧ�L�a�Q=�V�_v����������]�:ҩ'(N����ZX�1���Z }��!�ך=糖#ǙT�wɕ̿�b����7d�T�֪�T *�)�}DW�����W���������ôv,N��L��~�����
}d	�Ҷ�|�O���D�%�
Ʊ'�k��eV^|/D�S��?Q��g,��6`TE"��
� �.j�+��EZ��a	�m�V�nb+���3��F��|���ZZ�Dt]��W���F�E2�$�f)�ƾ�(<���@��b�ɖ��ي'�'��b��:1��z����BdE�0b�{Sy1�QXmU�n�?=?�s��ebǆ�1�LrB�\8=&4q~�2Y�0����|8�	wk���ZZ��g)^�yB�����p�ƃ�F�5���TM��/��w0G�����)�o'E''�s~0'^���P�I%&ƗE���nv�j�@+���y�N�
���,G���^3�3-����'��ѭ8�|��m/�|B<;H���! [D���ؗW�5;X��X,吵?fR��۾��e�?u_w(��^r��Kھ~@`�Թ�a��}dX1�df���7�oa�O_mE2$<?_����ls� ��QmF�r9��oJ<�=[.�٠�c���^��C��X0f���{W=x��Qj��mx��ֿ��)|���8�,�S5�͔�qw�y̸���q�N�]��ƼIkj�.j�������ܘ����� fN���������IPǋmK���w�l"�ahqq\�N:.�/�](s=�v{�|+���晄p=ػ�rig�Q�3-�[��L�r�����Q%��З�YŢ׈�"�R[*y��~��%.�.e�.�����d��"9���iXt�[F���4�0�8>����S����&�gz�r��ʗ������B�Hxbg�r�F����
uT�N�a���j�wҲ_� ՛6�.�g�_��ڑ���|�;DW��x� ����[��]R�s�%��l{��Z:�D0F�d3�Q�va]���Ty|S�4���˛�h��؃y���C�d7CF��H�tWs�h��o�m\C��ו�=�B�i�� �A��8����h4^�'�b̀�9?�Y�֯��7�xS��SI0�w�1d}�F�G$S4O�U.<�ZP��ȯ���!��+jq&�����PS5WN[@� J,����	��?��E�,�>�-+���,�X�i˟���с��:��5���m̩@2ZZ���DX����l�{�L�&M���h?�ۅ]ԣ��@>J�Y
��r�|Go ��vQ����S,7=��통����%j�7��b �j�.G"O�8�n�U{�R�q�c�(�[+�er�+{BW�f����������̘\�'k�x��2�����Y��P����C��-Z`�h'W�L"��.Q�XMW�P=s`4�NvM�mQ����
ǝ��/����m����N�/�|	G<]�{6�j���xW�3WS��T�[D�� cn�p�]++Ec�5��C�j�Ç"�^_F��a�{)���()žp��d���I8NG�#�`q���<��Φ�@RhF�<���h��4C�.��SdW��ț8�������Ra��O�<F�2�Z���OZ�3Y�x��~�z��:O������^���FF%%>��^�Q��#���d�ɮo�������MV]�R�[����;�Y�0�c�x�a����< �6w)ސ�z��D��RѬ��*�M&5��ߐ�k�*d"�]|��0rJryJC��W�¾��,~D�����+�eز��{>5<�W|��Fbj�vƌ.Ԅ6$����N�W�����l$▴�� ]OQ�F�|���Diᩧ�Պ�a����:��G�l̵�ܵ
���WJ9v�S�����ޫ�$��,��>��H1��E��5+�G�@�w�j������Ta�B�3�:,(���rD*�`�,��OPU�dmkm`����$;^dv��5�Q�:�#��9�)w�ў$%�s<_��i�V���$�C���0m�+*>���X`��}�5�l+����vL���U�Y!h�n[��n]/@qԣҪ3$ %4�N�3����&�ߑw�/Vi1.S��W;ղ�N�tumF�&h9	��$暣�ԟ�aX�Z�B��/�tC6�_��RQx:Sg����`h�V�K#W�"��v,d��*���<��1����2�(�\�M�N0��)��s�+�_H�D��4R���⑰pi�m.���l}CT��:�z�
Y�V!��tj<���nh���y�5:��T�zp�f�5o��y�~�:4b ���퐖�Լf��޷L̨H��A�Y"�
����t)����;49q�r��9ה#r�	kY~	��qW`F���C��"�wg���5��qQ�;���=ť-�Z��{ޚ� e�U+�
�>���a�c�Y�W���Yv��۫����l��îaT����O�L��� �u;h��jOst8nm���zm�ͻ�W�_��{��Gx�Ar�L:00����J�W���:{�,#w}R�>H��hf��ٻBgh�Q�G�^ycYJs ���;M���^n�:�oVy>��j��݊����]�F�D��$�����-J
��i??�ll�@4ω>�=�J3���B��+�F���T�N�7Zv���]�3U���L�e�M�j�k�	7��ɓ�R�;B	�����9�:p���Ua,W͒��F$53f��ݭY�Ûw��l}�k~f5���DE�~��0���l�R�Bx��,����I�8�~�oz_�nJ��P�>�7bn%��ܽ)��z�Y:��{�
���&�{���6W%0���L��oB�c��@)4�X�(Ϡ����¯�9����D��@��CG$�	�����Y��=�o��;�C��{���\ߓ	v#�Ɨ�@ٗ�{��ڟ�]�FOk��x�xx�� �6�� +�������R��%��k�ֹ�f����]ѳ��m��3͘���Y�v(��8��!��} �_|ˀnC��O߳2z���L@����p@���(W��F��4Y�z�P網��D��T,@� ���p/8�+�q	�u'
���M����	G�,�xz6E���D�.�7 �����KU����{��Ч&<��gk%�%H��.��ꗿ�+��L
̓bGT���*�O��p`��3��$�܀��]-Ԙ����}Z��������x���9	��fn�"��j%�Z|��I,�w'yz�M���h����t�vt}��&�c���f"�1V M�Q�}�z�l@]�SC�*f��7gI�Sn�F���Y�lƑ0.4E�GЀ��yM8�^�*���4!��c ~7�M�2�h�Y�m[���L��)G^�2�R��+��+ � ���v�vx���7��K�h��ܳ�8q��A�x�	�2��Lj��+�w��Ӭж�'&�݄S�{w�4�*��pě���rZ!.m?|i�&ob��M��@?[n⧷i�����������V�m%ܡ�^-�ڥ� ��LA�i�F�����4�n��Q��H{
EO�6G}����_'^�*�%�L�H4r>u<{�����<s�L,2��j�{� XR�
�;�}4S���K�Q���2)��O��woTxF��/u�k5��}��HA��/m���;��5�G�1u�؄��O�}�m�*��-B��%>QV�IM��'�ܧ�
e��s�%��4���jV
dԧ���u8�Vx����."|�j� }�Y\L� %�,�*&���U���[�!V9�!�*Q��8�ͼB�#��1R�$BIKS�kKDi,��D&�v��*;|�0z[��\���t���a����'�W��J}�\���e�I���u��̰J���W�"��'����C'��DCć����aA[^'g��[D���6�B�5:Y�����S�U����K�e�6f�%��-2�i�.�*;<@��)�"�s�{�K�A���t�ʚ8��[LO���U���^�Ŏ2 	�<��]��x!Ӷ}�:�8��@�4�x��6��>H �An�4 ��\��?��&xA$�7�=��M\*p��iڒ;�^}�O	Г��&.isPT�5Tb��3��s��󶆶�D؉G�k�q%�Ne����>��G��^�����$�kZ��������B8M1y�\�i$�0���>���=96AU�Gf�h.�m�-Z��K��dw�
4���U��՜��U��Q�|c���RL�hL���b~h�b�J9*�1N&���i�o�[�p4:Q�$$��Nk�2>�����7�H�o_�_+�}�B�k4?�Ϥ��s��}��9��%��1A�Dx'�J�%9���UK֦y�p�9 @�m򮠧�ϙ��Z`��b5�>Z�(w1��Z��+��)�@TZ,���)���Th�sj��+1	�?�%��%&"����Ej4��'�&5�m���Kv�d	[�d���[��-Xg(�^���.��Ʉ�\j�V�{��v����(�V��( ?*@�BZ���9�~��q�"��%��%�����T
��1��%�%$P_~�������(u+��Qit��W@ )��O�����������,_G�9����~ê�+aLQ���)P�������4-� ��B�9��#/���fՑs4- �!mF#������
N"��K�a9�j\�B��H����%z{f�n��oV ���fTL�Ș�:s�@ӷ�`%�>[1~ʻ��R�m�ɖf�����J�MVj�ɹG������V���^9z�mK�E�>��p��72����0R����
|ؽ@��ހE�p�#�īF�&pY�j����@igM����h�[�-��w����0Q%�"�1���lhE�;͋�-JDp�����P��F��kh�Q��@-+�5mO":��߳����Ω��`���A�:��5�ƽ��m����@@C�P�3o[���-�Ծ��ht&Б���U�@����3�J�joab�0���;��޽w����s�?��-)�Xƞ��Z���柌?J�y9�\Y;�v�u9[�Ѹh(�ԬNWa?�oj������{�O��w@�D��i�/�%ʽ�|#LCFM��"�}�+��aVA� <�p��J\��� ڛ��h�\���~�
Zh� H�?)����#��fM�K��RESt�7X�'�7鰶P��:�0r�[�Y��1^��1�:j��-��0~@�H똻�N��)����o��/_��������+�u��_
��e~}7<�xV��6|� `piT�J�h�<{ �^����U�I5*{=yմ�O3�څ�?j�NEh�|��wc��+kE��+���48���� �K�غB>g�'��z ��U����}���D�c����
k���%ga���Ev^��5V���B���(1��A����g��1y�%��So�Y�%M���ދ��ñ1�\�v<QD������~������{*J�[S��4� 7Ӷ���|�Ụ�����H�y�u+��tNI�O�d-m���%�;��?>
t@���ST(y=N`a�Q �����|	~�c*զ����֗N��;��BL�\�݁gј]�v�#ǳ��@0������`c���^�^�C&UJ�x��:�Y4f�wh��nҊ74�@�,߮���9�������s����} +������r���o�g��Ju㟑�;��^��ۧí���� }+mR�!�k�N:�r�ډ�f��-d�
�_�+Qߝ}B�߉��
1���N��W��S�\�.�S����擵Ϋ`�f���;�h�
,�'�.j�H�6H��I��Â@�
I�ߗ���^'�`M�6"�u'7V�yT� P��s|ՊG�9��qP��na^x���l:"�Qo�:u�T�+� ���K��ٯG�����}�u~3�Q������K#b�)�]RY?��=���7ˌ��6�C	�>�9��9�>k�7��$"�wў�\;�?��g���/�MMڕ�p?n�h�1<dd4�-���0�:�+\@b�W̙kXk�l��r;
d֤��AFfJ�\~YJ��i�*4Bpھ�i�0�����0��J@�e^e�қ̴WlmbCn��u)�\��4;`ծE1Ç�t>���	�_�Y �:�3������7��L����g�u��J�TD��o{@�9�:���/Wqe�{�. �l[lݳB���5�F�
�q|�4�:�iu
`8�>���=���XE��Q�yB��?�"�=B�j$r�ݮ�31��{&Ҋ��7��g]-$?�2�v��!�L��{��4M���ϴBsg`�i{��ɩ�B��l�������F,*9�jt�t��E.[T����]��u���(
�i�zI�=扰�?��!_���σ�bi���6���c�Np ]Y�<���@���!���Ȣ3/���ǧ@���*d���'
lh�0�0�p\k����S�V4S��6�[��8~W�-@Su�)�I$� �AG%���*��䗙9-9g��� ��B@��ep��S;w�� �˕*�)��*x��:)kī��c�Js��	h~�ƅ���|�<j�/.D@U���U`ż���n�W�"%�ζ_���?S�R����=i����j����`�g�)�ͧx�䓷�f�:[�yxy[�,֨�7�	k4�5M��,��r�_��a߉A��C��d/�S��b����Lr�a�(~j�c�v9��S �~C�4 �`����(��*-�A4w,6����H=,���i�`�F7�/��n���`3%��HOz�D8�~;ܪ����w����/P�h��EI��D4�;��g~w3,���(��Z��!�htR�"i�M�� OF1N,+�}�y�� ^����d8��&;��f�&$�=�8��S�@�Oa�?2Gi�Ki��5ؤ�S�5�Q|�ys��ZV���$-| .�S]�|n��%:B���-�W�����T�\ ���O�:�2�n�<U7���R���u��//��C���p��d��d8o�o��腂�iXsES�\
b;��j���F�Đi��v�s���,�d�U�U�(J�ҁ�h��GT��ȅ9a�U�9��7J�z�ZQ��'�`�T0�
�,�C�:G�kG�/�.��k@)S������@��P�kN�6L��J������X���A��9M�0�͗��S�L�����D�N��A�b\d�R_��SI�u���H�z�?PuM�}�gЃ�<��TF���2d:����]���3�)��|l�6t6[���n��I+S�W�Jk��|7�{��y���m���~j<����U�}�N"	%|篝ZI:Z�Օ/�P�`H)^��IW��s�.���DYW[܉��D[]���6�b�w��UYCF���j	p��a�����V��&�9eT�yη��_��7��/�	�3�@�3^����L��U/&���7h�8`�҉0J^��ӥ���hL �����*��T�;iF*r�N-I��r?@?����χ݋���N>I����ʼ�����3�:\����OU��χ]�!_3��FMS�
��+
�A�K2���=E�_��F �����<�"���h����q�G���+@����K^+0j�V�Ou�'�q^��& RM�@��+��|j	�	ȵCmxmie0w�
�G�*郥绖�5���rU�c�l'�t"X4 �XQ��x�x�5rv,�
jmeH9$��:@�=��E�)��h��E�P�QK�����<^����p� &�S��D�S/}><@/e,�f���Q}.mz���쌍�KK�^�&�uj	gnW�G}	�Ӛ�i�5W�ՇW����x{utS� ����;B��;�N�%7�ѼR������!O��bT������y!�Dr������\�-N	~:��4��ҨzOh���*2��8c
t@?��������iR���X
�}�a� ������4s���T��߶����
���1W! ��}�:�
&*@_|��}�w���v8�����&��oS[����__��Z>�@�K8/\M?�ʹ���̙���@'-ʭJ1�b���5���WYk�to�u-T�|��S��r��72����g�l!ǥL��8�0S��]#����r,oH�#ҝ�d:�ҹ\A�-Hl ��N�ܝ��4��Є24�/�lȐ�~[�`|A��>����2Z ���׊�)�mG@\݃B-���m�X�)͛�, ��*&�X=�U׳��R�ZD+Y8�����h���%���߼�`����e9`��E�:���1Q���u��2}�8�R��V�����ZV��B���-\[�X�v���)�Jm�d�m�e�V[7*��Nf<j"`L�7M�����?��7(b�_���������)������'�$L�[�� �`{j_G;KZL<ZY�Z�C@<������*V��|�ۮ{��-G�e/&�S��A�8"�o���3�
���̛3w�k�7��p)^�	����@s5ʸx%0.]9蘹U�Kf����oT�C>�b�1kt��񒓾{�|��2�.��F{V���7vǭt�%/�B8�&���ךq}�fX�x7���>}���{L�-�?̞�{|���BC'�98�$09��iL01�2���؂���b]�z�-� #)��)�K�aL��������^Bʼ�V��3�4�� r�h����{��*Td[in�w�i�)`	2��AS_�4��F���j�����ԽN����2�,��+����\���a�����J9�dL!��ϤҚ�2�{�`����v��Opۑnj��k�2�e����3��|�6@�^��5�l���$�8�Z�G������M(�P��)��c[�{�����)��g�����?����p��W�:>fG����esμ�Þx3Ӡ�B,����	@u'_���~?\�������+i��N��̭�/�{�n��u3T51h)�?�_=^&���0������/�����U��˼�f*_�a������1�3
T�Ѹ���T�
	҄đ����9nf���d@K�[��R���R�P��2�>�]�ݩA�p�	X���D�+�j'��J󿲽�:p�<�b|D����ʲ�4� V4'8
S����F�8��e1���T#��U��!�TiU��Dӡ����Vr/]�)����6��P&G;W��%\)2�K ۰��L�.�W�V�Z	g�@���|~3l����ľR{�[�.e\�̹�։���4t7*��!5�+GJB@Ŕ��4��ߩ8�8 |�X����6�%i�L���f��{����}҄d�<q	�V^>�,M�M�|��w������Xh�/r'���E�;:���
��*�8�y��i�����%������- ����=J���|x4��]�&*V,_�����D��۾0S�[y�}]��W�����S�})�~/ƚ�����W���/_�B�Τݽ|��9҆�%�Mie;E��B���&���d���˃M��ܦ��>F�ud���? >�´ь��v��e8��F��g�xW�͑���\/i�����!����*m�:� ���R;�n1+���v��G�J|b	X����Jm/�	�Z��)m�`�h���7��-��需�D��V�g��cP��lT|�=8@G���s�L6쯦�]m�޸��~>���%����s�[���%�N<�T�WZ�VibuL[�B���v[S2O�yV-.��� ��|�5��]��������U���-P�91Xl����@$~�tj--k,�w�Ⱦ/�G���=��b)��xp~��)b�~c��׿Sx��V�;:���
d~���1?�����k�v*vIV*�����h�"�4���3F��ћ	�{�|�䶆20Y�;�C�w�+��|�b,K��ԝ������寽P@�R�̭J�"hiu�r�=�	V)C��t/kN�Բt��j_*0Wm�L�GE���J'{�5R��+w]�|�ֺj�ݧ�Bj�w�{��B�[ �A~x�q�>����6w��t�1"�u͝r�W�����t>�S9QY�
��uW��hMn�E"��D��k��E�:�:�	W�a"��G������Y3k�-2k���S5���X�*3�y�ظR ��8[E�S3 ��1Hg�e���%�?�q�l���p������;����q��e��/���F�>�Z+吚 ��yb���o-�-$��>!K��v��-�B�} Gu�5H���}�֡5cR@��8��4�1�*w�[�.��,4����R{�
.Ҧ4B�	�_@��f�M�e-h����z�c��3�3|�I5���JK�	D �p�n�F��H��8s
t@?������sdB�D<���Y������:1��x+.Ѝ@�����5�O���Z�2����[�˿U��"��O�'��9-3��ff��.u�:\���"�
��?8l�u�Y��7o�0l����T'� ? #�)x+�M" �4~A��K��d�6h�.9�xk�\�C�<" �'EO������Z�ז���R�ZB����iWc�KH8RE�B�#�+��̓�;0l��ۏ]>qk��j��.���]�彗�-_	m��X�ճ��
�%eo�h�1�&8�i�H��-@']�fZ�g�i��((��(C��*�9N�Tp�L��qT��^��r�l�YJ��H@z�w=��Ϳ�_biQ�J�i\��Ĥ �Tu�L]���>w�3�R���XzZ9a�Z �#�?O4{*:n�)�M6yE�p;�y[Ĭ	��_�%_)����~*M0h�55˷kx�E@��ײ~�i�SV��HX(��r_u@���\_v@?ו��ya��K ���b�D������	�B����v�=��"#r �\ReY�2�S�k�4.��w�`v+���v�iF���+mOҢ�߹|����代B�?� ZAp��[�d=|��a���*�'��
����Ю�%N��̤�/��6�2-���욣[�Zs#��� ��Al�|�t�z~5�d��O�y	3	
i�!S.>^kqQ�x�(���m�w=M+xͩc^���Nֻ <��x���7A��3荘�ɶ��5/	#-
ݑӨz�����Etx�{ېx �Z߫?�3YQS�0��Ạ��r��ӖT���+�qO'3��B��߾v����o����vx�=�&-Z�']��B�$�7�"DTL�[�x*��SO�w�s]	:R��FMw�Bx�MB�kY��@XQl�H�&Ϛv��Bo�T�� ZO/��B�h����]i��5{���=P¥/S�
?	/��p帺�R�����'��W}��e%�<�@�0��84e�i8'|�G
0Ta���\�IД۞:�9҅H��
�#�I*�j���)XmM�8��m�y'0�[}/���W�x�k�AZ��r���t��_5�ʹ�|���)=M%9o��o��OЮ�Hw��q. �ħ*�ړSN_u��:�A�E����̹ҮŐ��3AO��Ŗ��(���Ӎ_U��꼥 .��/���ox�L�b�O��2d&�Е:��h���6Gė�����V�04W�S�/�em�Z���5�"��1-a�hfi� f�S��"6�
�H��8{����|�u%ߝ�?�ۦH�s�m��T��K�I�5��R�����h~��ۿV����\k�l#�w��,8�x赗brF�+B���&�#�GN=�j��]_9&x�� �1�b:U ��������������8���b��7p�#Ƽ���2_.�XTh��I���y!���Q2�τ��d!�4�H�B ��h�6������W�#/�"��a��'̌�A���Ct����S#���\=�
�[��ҁ���O�+�}x�bX�O�z���I-|ޗ��:��׎d��$��Fy��;W���6���J�E� σ��#l4G)W�g�:�h��B F�9�U�K�9�_�i�?:���t�ҩ"��<~�����/d]P��4S�k���&�)k�`^0u�?�o�V��G++
U�bZ��1���Oik�����8�C�0��jM��E���#�������"� �{� T�!K��ɽ�WZ������H(m��8����0_�:�6Z�������W9̿�j�V�".�KL�T���C�@E�S�����&�V�@������`���0��lΣ#�^������;���D��W�j@GH-�7Y�dL��cH8w�>\�����|��f���dP�����JXh�߻RL�y:W���D��<���s��A�v��G>� �ݲeI6���-_:j�� 844)��F4� �A�8F�����~�K��v��]D���X�v���o����0���/�Ƥ����Ϭ��EsG.]K)`�b���VAS_~3<���T�Ns=�B�L!�;cǼJǴ�� F�o���׊T�@�c��aWJ8���WZ����3D"�X[H� e�6��r�x���v�}x��~U�#j��.��ͮ��Z  �vY#,�j&)�2o�����>Ƹ >���;�U�H�Ӫ	yV��`���������`m U�4�N�;.	=�&�H�m��. K����{�%�4�@�A���@ ���H�Y�^�j���������.��/�ƈ�>��Zrp����H*RYo�kbA8����,�\ g�V�D��7��l�����K�q_R8G��/�����{�Y�j��!.�]�.\7��s�ݴ6�ɣ�j/]��~���܇��������XEX<�\�+j/}\2����/n��s[�?�x�e��fxA��]����-a��@�n��X��ӆ%N��E�~O>���e��%L\x%f�J.�B1zS�r�T�E	K��İވ�_�l�J��d�=ȷz)��� ���Z�Ջ����}%����*��	�לfT�-ifT�s�.�ҥi.����:�FO�ߕ�pT����`�u�8s_��h����"��#pEC�lx�T�����a��Z��ůک�w���v�z�k��CW����0r��R��~<�~��55Õk?����I�*?m���9�f�".T�k�[�[�󚳮�v�����Q��/ڢ�/
ts��L��l�}��@���B�T�˜������b�q{Br�ܿ�ʨ�c{�N����+�U�,s��_�5�V��'��*h����2�+�ʹJ`��{�6����i�*J�1���#���#�$D̕;��""k΅�����<��^�9���? �pĚ#�a��%��;gF&�Y�
�����9�c��	�l��<4���Y���;Dz���&J:�tGю�N7Rt�b:��	x�?�Kt@�ǾB�6�'@׏_J�����9ٵ�Ø̎ ��/������2��)�xbVu�,ik�S��߇��v�s1"�C�������+F�R���;iq��'�n����j�7W{<)�v% ]I��Mɉ�����B��[]_�o	�\��!--�Ǜc�(2bWWv$4�ݐ�#�&�0��27J��ҡ�1j�,�8��	+MaÅL0I׺�����|a7¨V���=�t�	D.(���ʆ$�b�ד�q	N��)�C1��Ŵ�0��,�|#k����/���������2k������
ܚ�p��[.�w7�����vFE�K�.���K�.���I��0#K8��[={��[U�{jm�������������E���Xof��KxS��2(��/v7�l�A�e���e�57!�ՑM^�]V+@�vuc�\?�2���`-ٶ����5>���f+�/�G0�����������C�s���9�揜KE�.��M�%ŐF�^i�x�	��s���'P/ yO1e�k ����P`D�,�])XBʯbE��w��Nmm�'�jMn3EE\�EWTԻӢ(�t)[
��.4�B��c�(�MT�h�	�R�Ա �v��_X(��]T$��(e��?�gӭ��=��UN�',߻z8ҙ /sr�@�Np6�
d����hd�=@��������0M�;;β����,���'�#�hF�3n=��}� ��F�*��TOq��l�8GH��H���zҰ���v�7_~i����S	jGYb0sK�����Ff ��lBf`�5�S��JA�[�Ln~���J�ӵ�E�A֑�\1k	$��w�^w����d��뿓eG�+ɭ�|�ͷ.
���h��:r�2c�FFh:�<����-0>B{�֤��Q,C�6R#�����)rvGR�,�>D �x�c���&��9R��9���3�(�8�)癟|�Hc0���3m����	�▉�.c�D۰i��3�H����JY��M��1c���Oc]ܪ(�-�e�(�F�%Z2��:z�U�̚,xh���A	r�=U�#�=~�\� �ƳF�7�%b�>Xk���b�  �K�Z��)N	u9�����<`�ָ��-��)�"-�Z�l�_�s�T|"b^k � 4}-9�Ρ� ���5�'�;���^��C֒6�YO|�c/z�)`�Ҳt-�H˥	K��vҕ�n%-}%�\]����y��4�2�/U�r��Z�BY)z��@,�r���{"&�t������0����ߪv��I*�J��K7�N�u�Cѐһ*8�VB�ut�>����seʚQE}��Y�$��b�)ߣ���+��#n��c�jk��#�0��{�
�?���@�8�}�o�o{�Xߪr��?Κ��zy�ora �����SFcp(0t�2��I1�('��p^����$˄9
pR� fC�(͔��v/1��su:>V��M�Ơ��]��y܀>t��=f� Cx`��a9�̾T�����9W�A cpX�cn�s������csj�����~\��F�U���'��mb�癴+�V-*ǲ0BqtD��}^[#��y]�Ю�_���z��I��t)[���iP�ro���� ��"�A�S\�����_/d_*�`qxg��N�T�R��򯩺��V��K�x�f-����]�'�hBc��)+����T9�аW����"�I a$���<h�/p+�w�BBg�Xblm���mz:�]T��S���ٮ~��QCo�o@=Ҝ�_򧄇��hN��>d+�>a]M���4/�U��<>v����P���,�O�,+))�Z����z�Fm`
��"Sk�?=f
��6�a[#����O��H�Vf C+���!���}�4s:��6?<�oG3$Z_1;n� �k�C۔V~��wڸWW��V�[3������9�L�|�� �A�"�6ۂ��ܖ� 
��
���'_��̟u�rESox� ��j�7�qαe�����f�ik?=��X#e!`ng�D����яyrQ�e-�zXE���zBu<��a:�̦��;u��2o�2�Ca�/��mD2�	�4���>ۉn���N�U�Hm�#r���BA��u:W�!�O�{���o���1V�uh./K\I������[�=ժ�n���	cm�k8���;s���Ҹk������]9�\?�&GR)+�w���riW�=��?>#
t@?����S�I���e
7�/Fs2���-�֠b���O��������s/�i
����\�]\Ӛ�s��.AP;������U��y^Et�3<��� ��������{�8����x[Й9�N��^9�vN�U�@�5�l*H��!������@�h�o��� ˚���)\C.@�W�b1�6��i7�E�@���d������]K?�{��)|l�f��`�\���F��J�h6h��V����t'�s�2;��O>�
4�S��Z��r;嗓z���vF׼����>�w�+"�r�*�(Z��K� 7���3W�J�K�`N�r�I{��-�Mp���f�J����[@lb�c�T�Ю�X��Tz�o�^�ym�� Ei呣ʬ�IF��Q9U��>�ᙾ�~���ӊ��x1�0�Ɓ�ݴ��^s¬���A�T�]=Ph-���)PK�N���ё9��IsW:���k�3��^>�񔆞ЦF���QC���lL0ۃZ{���������W�{�xi���箕����i����fL𛁫�t�n��G��iwm1�Y��M��4�,B���;��@�#��N�E�
���Z��p��dl(ժ;ю��}0ϳ��ަj�H�S��A����Sq���rs�jvy�ua�&q*�fA��*2�p�P��!���XL(�-�{&���l��]�ᡕ˹��tL�-k/���&��c���+	*N�u*H}�8�]�ju��f�SԔ�q��x����K���u��:��ݒ��	9F7('5�cb|K��?ШU 6��J��n�`���~�O�3cG;2L�)�iAQIq���2�_�&����*�l���L�NM�I�2���V'g����
��`�5�%&r�ў��Y��.�M�������`q@53�U.r�˾p[&P������- �Fs��������9�r��������Wj��J�6�&��At����ؒ��9�kܷ��2�F>�������\"�SW]�Q����3�; k:V�&��Vw\�P���Z= �W�9�
9�=�-��� LZ�J�0��s�e�J����� �P��E�����sӾ~�]=��>���L-�q���ଗ7z���V��7.��0���m}]��:��c��p\��F�?;
t@?���)�� �=�����A���ʒ ��{����$24-��wrL����Y�m��ET88 ��ּƧE4����@kFY"��k�+�d�0�b������G:�?�t\ 5����ј�_8�Nf���'�1��$Lրhm8љAw}��վ����R�y�_ ��.aSO�A���)|em@ qz`k��1��3��D�����hB	]�.s�?�d���#&|4�5.��D�+^�8�% gA�A�&��#��0S����ؼN��HC��V�f5������4d� ��qyԢk���"����@������8��	�Y��O��7�M�cِ��@-��-���f�ɍ�U���8{
t@?�%�^  %b��4?���ݘ���Y�w!j1| ������ɴEE����}��y�_�sR _x��F��/��a>\s�h���Sװ�k�@k���A���ͣ����m�#��ĜL��1��V�Â�T��)0	F`r���.8W��(:�Z_�����:����$4�t�Q^�&��8�t��<�`a�L�m=#d���U�̢����U�ϸ��@��r٭}������{����CK�Z��-�[��!D�$�a 4��!����t�����-g�?���+�.{���=��?��F:�6�[�7�t�=���M$��[�AV���uƾ�*�8�%H�58����y:��_j[���+�\瓵�X�v=�}�k;ۗ��vi�b$���R�[ Z����J�%`�a��p:�nfW���u� �b���a��W�yiȅ�a�dWR��(�dq~���`0Ͱ���z��a����k��y\# k~o K��Y��'~�}�+R��~�)��K��Ӊ�ZuY�d1�!������4 �)�����L�aR}� k�v���r����<H�>j[8l���FW	V�.�´�ŏI[p�@��,gS��Z�v�Ghi��N)i�%�گ�m�V�$�=��X�݄���7i�����,�����]�-�*%h�ro*o�����nYe�����?� `��A��ɭ/̦`Q��v_��X~-_�1X,�O��G��+z��'O݂XB�l��D�I�����Vcq���\_��.^�"Tj/p�Ԗ�U#E���S���/�w'�	�Ѱa��W���CnsA4T�-y���ɟ*�a��{���zM�W:�� ec.�w[�8U?r��fud�c0�����cS�G<j5#��:(B�߇��o�3��6��?��f��/3�ڜ<e��� D�s.:ǹ�Zqi�v��	PDl;;)clͱ#(��e��}0�K� �"���:^�T��S��{"�OjF\�ހ���A32��#���t7g�+�^P�_�jdD
r����\�4MS>��0��ܖ��=;�wM �[��I����F.m�@:���Mj�$M�Z��4K0�EKc)�@�P�ⵉU�¡cr��p�f��Dz���j?� �J��ޏ��
"Mm{��[�ǒOY�bqP�Nl�!�gH��g���P'�6�[^M���H�*��Y5�4xX@eD䘀���$*ߘ��n�ATM����$��ӄ��ךŠ4QG��xNe3K����$��O���0�p�����c&ۢ�͈�)��hN�Z�y�@��o|fХ�Y�bbu]nS�}�Ԍ��R�c��(ksx��mQ�
�n�`�{`Tp��7�`� T�0� ���c��F`y֍R�^"��O�Wj�7�!�!E/2T@����Y x�\,�h�_Z���V z��M�����K`�6V��"� �,DX���ҌM�3c�k|�p�4�7�a
��f��;�v�`��ɡ�8O�}]���`�ҼC#b��os_���%�\�4�{*`O��òo,̙�u��7.e�֨E��"��YQ��Y-珛��BK�MZ\�M����x�_J��1�M�S����l�Pc:̈́'m�	s�>w��|�4�Lܚ\���)	�_��aVM�0V�ߖ��ϱt�z}?�����G�ӻ>B>��>9�� �(�d����R�4�*틱�t�jsq)@=ɋ��
赭:^Q�v�0@}����r��]h���2;���7�B�kY�t��Ӻ�󼁿@��0F�ۄ��`�����r�� �����G`s�EZݺ��P)[��� Y�hZ�v:,�~|J�Ø��]`����0e�,A�����-�O����،^��U�t�U�lZ��?���ner������<�x��d�m3>"F>�Oa�~��}/@�,�gM��g�������{��?�O�+�F�8K��*r��;a�@3ҁ��T�3�b�S��A�����O�}l�.���2Xhuy��&ҿZTp�~4��8��������0�ގ9K+t�8�������1-[�[��S��	|�*��X3��H�HD�WZ,:3�w���!���;�}��ww��Kp��{߹k�wC��]]U��I�M��a䌐:4I��a��L_�8��ۙ�Z�����B��P�H�GėrH�)J����v����㼷#�P��-����M��(��(Ip�lˌ��2b�;�A��D����p�|-H5Ʊ�s^�+�n7��ٸ�ï��^��L����X�*�6�U�f��c/uVm��u�>3�R��'Msz�L�y��n�[�q�
�T�c�X���9�&�&�7���tkK�A�����3гG	2�	}I�x{��O��`�W�v��4�Y�60���>"�v�M^�R��c�;1�&5�)G��R���ɀ�N�CTE� ��t=�g���sq��W}��#6�"ȵ���Kb�q�ެs��@�bn�&8����E.�g�k5�"���MkN�͆;���NX[� 1��2sf6�˞��+4PR���K��O�C&`��I+�9�%2c g �uYe*�Z�+�4�x���2��f����0�}��#Un:�R��a,���� �:��\G���v���J��V����?`s#�w�T��?�	�oZ�!JkY����ӂ�)F��Vc>A��,Y&�Β�2�t�h�����z[	 rX
Ehk�a�@G��d�C��A�"[�Nو�I�ԑ~֗:l�8/��Z4|`|j��Ɨ���)�z?'�{��~��߉�l�[�Ƀ�w�ξ�V�ۭ_�E=�����o�Z��f��T�3y����F��m�Zn\>�!�R1�m�%�]%p��-�:�����Jg-H�W�/�����|�����2�y�A��f��Y�a���@�7pw��)`���]R�L��}�!�̪���$<2H��\��ŚD�'��?���O�u4a6_�rN� ������u�3Fy��^��
�Gv�T��9��'�KG8��5<�Lf{ʽ�%b����pv�f���4�ƻ���⅕�o�r�����z}[�O���H? pM����­�^��x�0�c2Fbɾ=���yʙ>$�Dr�4^a�Ѧ~�4"ɕ���5��[s6��0�G4��8.�-O��N��3��Tp�D�N��k'E_mYEwљ[�c��09�~7�&����iKr����X���ڻ]'�ِ6���������1J��Y=�ߵ��Ֆo���7.?�c��m�����y�?,���,&��J���_j��F�"�ت-��\�ެ���W�N�$�� �9���yk���ۖ=��ĵ !f"�D�I<:8���#(_��HP�mֳ������i; F�%�=e`�fҠ�OE�F�C�!&~%� ]Wa��3p����2���8�]���\����m�D>��a���(��A<��Y��D�#�e�(b�[Q-]���B0�|����PS�1�F ����Up>��ʜ�ڦR-v��[;��C%�/�2�{�}�^\̡<�Jk��.�����|"#�&wq���W��/l���+D�i���	�+Sh�s�wnn��*�!K/U�� ���t�mH<���]��Ը��C̄������卭�Y���~&�^�j"vD��H�?��/�Ozr*��r�:���iD���6�:�9mm��J�W���#c-���GK$�Z��@�훅F1r7�޽G[�8��)/J`L��������{��~,M<�����:1��
�W�]^J��f������XiװU7�n$@-��uM�%ϻ��~؝���!�d�BAr�9�>#S.Juܜa��ĺ��{���9�̜ޅW5�	���t�e��)��W�d�����(��2AE����)�(��V�o��>Ôld���*����i��_��ݶ�1:guB� R{(�_r��KE� ٴ��F
��:�Z�{�]8u�ו��į�v�peIK�e���W.�M�Fb�.k��]w��M�P�3%|A���!y,y��MH!�,�����3MH����X�FR�3����L�/8�a5R��"^h�<�G��@b=����R$���p�,9�Y��؄��Ask�%R:T�Ё2�ȂMHF�i��)k6SP�ٖ4����zᝆ���� ��'3ު�yl����o�[)�,4�S�Y�+�;�\�g�ߐPO��9�����x����p�Mg�� �����TV�����.E��R×����.�;"{?ڻ0���E��n��R��1�2R��%u�Z$H�Jr��K���r�C��d)�ķO��TgN��z��'�����vu�$QڊA(����Q:�n*�9z%����Ir�EDL7X����%�{x�dsZ
��f�@<Sv��R	!3ک�C���2��w:C�8,	T�S$�aܬQl� R0��Δj6��-vf���Ǖ�(��i����*Ô#���i�g�'"���>���d�*�Z�=�c)	Q��:�a�uJ������R�Dk��l������� �lh���S����@��~�� E����!����k�q?T���i_zu��36��^G��Q@�G�>BD�0���0Q8��_r�shw+ "��4'6�k�<Ę�h�Ou��S��>*��:CԸ��C��։8�Q4��1}X`_�&��>�T�c�������mq��7��6�o�m���Wi�n^h��������7%�Ԁ`���g<T��ZX���m{Y#�o�>m����J���}r�x�����6%xyrs�	�b��,�D���t��Q��I�Q=���s#�3)�j&IەGrfUW�Z���=�-�6s��/N%o�щ�^��6� LCI�����q�K��%㽐���9��,^��CeM������	���<%��ʕ�F�?^RC�	�.���2�d�:�R�m�f�4���
I f95��7�W�L�+J�'\z�߂Ƥ-:̗�б�1�<@n���}��![�_��e`�uC�%�z40J��k��U��H�%a9����m�/m ݗ� b��%��	h���}vV�
�|��n&�JB�����W�F���X�kY�L��G��JP���&o2nU���UL���N]×)�_����t���<�K����U�����w����=ilw0A[���n�{���L^_>>t>�>�jyo��z^2�����ε�=�J�q)�f����O�4N�Q��nq��'�1�(Q�G?�n7���*ZϏ:H��q��pwJU0��� `�[ZI$��Q��ʻ���p���N��X��s�Ǉׂ���n�Bi>M�P;����N���r[)��pv/WdW�N�|��|�Օ�lKwmG�$���3������3Ϧ8V�7{�tQ����Kz8���щ#"�"ŀ���\�*~p(ׁB`�8K�V �	�ށ4�iKg���\������X�Q�Hƺ8J
��|8��D�^��qʺ�H��7�:HV���Ү
����\a���9YN�e:��	D��_�4K s��v��M|qˇ�.ӟ%�x��0��;�Ѳ;�� T�Y~Y���/3F���}�OM�x=?�(Ef#��R�#�l�D�~��/�dU������n�Š��� ��=����i(a����q�!�뗅u�ڞ ݚn\��F\���01G���^)�6:Se���A���p��؝eN��bG���ϻ�L��(!�����-�W�jG(! ���ik�_K�93�y{.ֿ�E�3�m�Fʨ��H�%�����̟[d�����|M�@$�����9���A�ֳ�\�ʝы�:�_���/�c�S~ Z���ÑUurR�\�%���翜������|9\.�+�I�׵�B�6�Ѭ�d�� �X4���J�M��IY!�8�I�kbJ�U닇�햇�׳M�.�Y<��orI�>8p��I��i4L�]��2�]�#F`]�P�/TV���純���+׊c��d�-lH�D�`C/5e��x$Z�&��!��T�+�$�Şf�`�p�����ѕ?�r0֙ta��s�ǏƜ�Y�/��{���:>/�hƗ�'� �qu��5�3*O���J\��k�Eb�b{����kR��B�i�彩g�� #�_Z���c֩C�-1�h��{*�� E��^K<Ae�oS&�$�,��M7�$�W�ں��d��>r7�"�xl�,oe՜�L�|/��5���J>fTH�a�T�u:�V���i�h=U	$?/MU6�*d���3������Ŧ�)�TN�q�_�EbY�}�*�u��Q��-Du��������F���2	p�#�W��5��č��?�|@ʵJ���bD��VK\ޑ�E�Tv���~��/5��}�(]&£!&�v;�-eN���ytW���F�u��ܒ	S�UY��j�X`���� c��Ϝ��>_==}�,�{(���Bt/�%*<�xf�%<��]�M��l�\�_���J��Z�i��a����]#��LMC6�T��BKB4��d�W���1eii�M-*�r ���>�|�З�=���_��3VܻN����8oj�~�_��ǚ���:�>��,u�\{_�?�?U��)�9bd1�{7���ح�v����s������ޭ��*b��tp�u����x�Ovf���ᷛ�9� l��L�����>R��) ��K�pd>n~L0�4B�7Rb����Ģ�Zz+����EY˅�'2N�1�|����O��^��������@�C���OL��5"�d�5��dw2�Br��	��dGFG!E��/�_��6ͧL��w,���n�H#L�Yʝ/�@�e��2��}�&PꍊP�L�i3����P���a����q��l���Tx
�_pˡ`y��?�N���`�:䞭������R`�6y	L�C�rn�]C�4֦V��3��B�]c^E%��H��-��\�J�drᨣ�v�
�t��辣�A��ϭ�"�1��E���ꨚ��+�A�5�	���u �%�>'/��;����Q_v���+�HO�P�xr�9��&���:��Q(4��[���}������7�4�d���m`d���2�1cf���_�!݄���u�/ȟ�0ce�8Iw��܁��l7�����"�2`�d�5/�8�A��� _5^;��|I� ��(�Wb�3�;�ٰ(E4��Mҳ��"I��π��+�W��\t��i��֢{$�+`�C��z��p�L&�©�Ԃ������zn~��������3~�ϐ!s�3Q���ZkJ��.��m�3O�⬱���~WOY�"�.<n�,��4�Ŕx�^��,�8�F�k~�Ɓ�����WI�F�'���el�=OO�.�6wq�9�3�2&Kק��$����]_+�ۜC%�+�������VrH��7��q�y����c�1_>x�nM�%�������-8^�e���،�5s.��]	W��oE���FԮ J�&\�ab��Z3b0B���3��V[k)��%?R�t|��/�ރ��*��Q�q|�6`&Kv��)�[�M�n���$R���[�|� �R�gIJ淫g�(A��4렉μ)�?��d�|�ǵ	�QD�(���s�Bko��l�yB��Fh'��f�:�[&@�nt��Aʩ���L����)G�"���:�%?/�z$�;�EQ \���F���x�J�5�  E�>(J��ćQ|r�W�kJq�F�'��u�5�<^q��5n,	�^� �c�=��G��V�I��� R��|��횄��P��4�D�б���}��e��{_Ra��qD�g<"a>���_k>��3��<�i��.s*~�C8U�d��u���e�C�����7*���B_\�u�*ķ��X�J�t}��{�0Ҡ�d�G��85`�f�hoF��0�0P@�JmT�%1��a�~�3�I&�W*���?^��o�����)�<�y�ĸ��p5����Ig��Ԓ=�&��/�����c?E��V'�����Xҧ�C9��y��E[��dB��5��ث?����K�����({5>A��%�����F�� �WS�s%�MՍ��u����L�5>��Fi���$��F�1���;\ j����!��ӶA�?A$��X���A�N���i�E�M�*�pxu�*�|7gO�7�0~�v;�j@�2}X����E�_[��,��<��k���("O*�"�==��w�
C�U�n��h(&%S���ni�͸ 6y�v�֖])�w۩����z���N��TV?�q� .��0�_����[�1L�CY-���QN`	J�w�������&a���� �Yۤ��������:H�x����~�,K���6�ovX%c���#h}ٜ������{#+ս<,��-~/�J!᪘=*�9�f��4����z�)�F�P�æ<���?}Ǵ3u�~$Y�S�'�@��a �󌀹r��)�ggG�`�����{��S���F���iQN3��$�2)�>��g��\b:��2����`՟S�A�5�⽾�M�E�C���0���
cv�^�3OF 5 ��cY�� �c��G�EL�eL�0ss�Tz�����F���D�#�ZfJ���ɹMx{�AF�s3��6!D�C�ٸ˶�zą�TLdf�G�g��k��Ț�UHj`A/e؉$�W�WVy�J��
��]���e���o^��6�R��%��c��Q�x�!��t��'��Y<>�`@��|12zD��O��֮���i�0��*w�IW�ג�c��ܟ:�Wld�G|��.�ZDI��#�(�������W�)e�zL>Ɛ�q��Tl�y��`�W�%�j�N����W",=��Cp���n	9�I{�"�-�N�W�7�lf�z_'z:R���CP��As���J[�߆�v�ت07kw�$��[y1�p����O�_���!&.��,ӤMu�i���;[��Nq2�JU�ܤ�5��<���;n0�T6ۗ�a�YJ`�������]1�!���m.XkT�nG�e�R�T�E�I�
��a0�³�Q;!՚ٸ; 9b�޾�0D���d|����M?��u`eR�Wp��k�\6O@���\�?$Rҕ�fw��p��E_^�)��`�%�*����r�_&Ak�64��YHS0huH�J��F
��1���ީ������|k�r��Oo�v��{�XR?0���Q���a�6�´>a��D��Ԙ������  �W�9V~މjۂy�f���Rj��>^l��V������*$G�Cw?.e��4ѫ>p�ƭ�Z�G�6�䪂Ym	�d�qz3��7�fwbp�GL���:�'�f��s'!�k).l6q��y�/�%Ѵ��(q�!�{4�^�j�:~����{�Wh�\��,��ZnyU���uh�Km�̑�Ajn��d�%?�����ӒSy��\;'�@��(���)H
g�i�%���/>/�6����������r]̏=���.��d�*�bHĜ�i�D�D}���dY��������	Q�iէI^iS-SbUE�+)^�T�@{�o��.�����=�-�W�\ѽ4?�_�K�|�
�"�������'��K"�|/3c�����|>�q!��3�i�(O0��[Fa[�8������.evk��2��#kO�����ZJP���&4)����ެ���c����Z{�p�a��vÁq���3G�� j����am�w7%H$;6��n��LĽL{��]�(f~�������W�|�)?	H:;�N�����[�cq�\ow����dL�E�[<ϣZ٨�#K��kԷIp���qbj���W��)��q�
��?4@�Uu>��ڭ)9!Ҫ�9��3�ݩ��={p�K����QM`�ɱGG@;��ɑ���ұX;�h �Ն�r���N�~k���0�SW��u��oA�[��Z�D�ܰ�u����<Ğ4l�<[^�6�_>��x�oS�F�iԎ���'���?��y}?{Mh�8~�yBiv�û������UJي̺�QA8nK�ao;�@g��¹Vn�X�Y4`c�a�Pݮ�����،�>t��4��	Wܵ,ڗ��]Ƴ����odYZUU�x�S�T���E>jm�n��|��L�SMCWA躒�Pp��ϳ�wB4�&����S�.�T�EBC>��c6� �� �=�wX�3������Mew�:a�t���~в�B���y���Rx�#�� !�Jՙ���X���"I�������Lm0'�NwM]�f������,�#��]�A������q��&7�I-2� �'�%�R������R#]��J��IF�fVQ0p�t8p^D���Z~�g*�&�����e5[�0S�qZ=�O��'����L|��,:Op/�_7r7�C�ѳw��lo�W���Qզ�=$a�LT�A�Y�k^�s����X�r���A[3�_�Щ�=~TlR�(�ME ��\~�����d�$?7`�r�,�V.C��ó�jL�Vw&��95�~����_1͟�����L�����,pBK(��g?7����	���� 9y��@4
$,�Y��ŕ��.o�@b<Y޳[B��39��=G�][�L*���z��a�-����4�.���Ȁw\ov�<�:��2Ў	+�o:Z�kȴ^{#�j���xPc-d}t��*f���*��e�7���7A!���T�
(�h@і���v��L�-�����[� @j�>���Y�o��8�er<E�o_غ��i*�&��KވyX��v2m��<i�(t��Y�_�@�Ų<v!����82�����,X�����b���9����IvrA�и��_�pcK+ش��f�]���ɉ�*�����Z���ݟ����<��'b�i��'ud�0i�C����?�(m���..
�yQ��(�Xh��p���f�B��z�.w�7?@�AF�c�pFA��f;�4X�"���(Sz����J�@�вY`El�:�hً mi�_�$�P+���9���t�zȳ��@��o�ÜG�������0w��W������>�� '�'�)�N�OP������.����^G����z,4)�y�u�z����K����C�+��o��*�U�Q����	�����;}oU���y��?kI���x"�F��{�h�8�/���#�n#���dm4�S[tVCZ�M�I��4��2��@�N�͛XL�6ؒy������s�"2:Q���B��]��5bO��IQ3�p�{&b��^owc=j37��,'!ZoF��O�y�Vmj�7(��i�;T�'��ФsOm���Lo��"3�Ә�v���P�)M��h����2M��)!n��T��7�}F�,�j]4��.�����)%�w�M�Y��.�x|'��J���}�����ߚ��Κ��5] ��Ib�n�!!�X��O�.�`;a�K?��g���mq #^e̻_F:T�̫�4p�&e���˽f2'4W8�2{����8t���,<�ɛ����ŭ���pw�?$.��8bZ8� z�y Q5)����H���V�	%���D*���-�eF�f�Ɲ=h����e���3l����H�:��Ͽ*�A�ח.Y���^BDoD󶩗>�����W��Lvȹ�V��z:�g��b>~���-�8�w���v?9��b�!�`'����z$���u_��V�0��n��\*�T��F�(�V�����¢0�?�1f(�.)�s�;�M���<�T0F��^�����ݿI���0�� {2�']1�ǰ�N[�9�B�8E�瑴l]�|"�g[0n]S�*P�L�"g�ua��#'�>���?˚�^��],�h�At"'��2w !ìq�85�@(�y��5��ܡ2�ِ�gO�>�:I����2!WF�@:%��Pk��宨�(栋O����ey����N��|U�=h=O��hVA�]vm0ō�|�c��p��A�Aܖ��gɛ�o�A�迌�i�tPC`(yi���s�o=���ڈ�����&b��l��?�T"�ͅ]�//`��ӳ�q �W"�g�L�5m����v�H<�` #Q�r7�{l��Ō�VM�Q�T�b���۟�9����:m�
�������	����Z}y�x�pny�6�t`<&�K��j��P,��*�ġ��5Q �N��~Y*��&=�^�����w*�z����,��N��B�����z�X�⊆}}r-�b�֕V��*�i 5���[�G2O?%�b�>����@�{!���n�J�N%�F\UQ(q�}��� Sˬf�]�,(
�|�_;��^6�ys�
��&���4�y.3
J�t��$n���T���?wo�L�|"������纃o�W�;n��3�L����̕ώf���<�\��>�m�dlol�n��$y?��Ch�qR��C/`a�\����W�F	�W��XJ��^���|8.>O�%ֈ��fs��N���-����&8��������dHw)�,a��O��By;����Ɵ����) �����T��u:���GS�bO�L���xH8F��|l�q5NҒ߲}kӯlK ޘե-jH�^ri��8�,��hDkQ�d����`ٸ1]�E�X�~��G���pB��	Ե��oZ�^��c�\% ��1n��7�N��1񲓙�,	�,������Q�z]����b�ÿQ1��Y�����̑�뿝�T���G:�A�%σ��}������ٸ�b0�}V@�<�Cil(�|�{���R<�Q��M��v�y��zP'c��R%9'�Om.���I����h�Ȏe��B�}|P��L*�T�	g$���a}�m S��I�s"t(�:�a�l��u�ڮLM�h�c;�*���)P��Ê�"��唒:��ҵ����|�hr?G�����#b;,�&�K��pO(Ƴ��Ž�������;�?�`��j�g���s�+g�.�n"z��\�AH�܄��ᘻJ�m�$�l��H�)~�����+�d��*r����:��c	s4H���Udm��7 �PK46���ެzF�v�_��~<`��X ��6u�6<I�#]�������{ڼDj���
ȩ�+�k��݌�`�y�L�m���dp�����PM�/�g�K������,U��oN���������jv�ɳ�|f�n-�I�-
/�t�H͗�>�5��k���*�M���`p+c���o������bA��H�G@S�G\:���Ϗ�|53�<
 �J�����O��74X=�JQGF%��ś�Ϝk������j�L;������,�L#X��?g��,C�D��<�M����4��%��6�d,{)�s�ӷ���>�>�^���UĶ x�	�YG��A�3�����ߵ΁T@o�W�98E����y�-/���_�Ѕ���]i�ށ�+[�����5DW�
�:k� ��qQ7>�e���2�]��7���;zGG��c�_	��vC���+㏧��z,����%�t�m�$X�O2^���+�=��[��n�cK������c���Q����0����8���<RhZ���������u��^A�/H�/ט-\|�ۊ=<��͇�uتy�H4�������ih�p�Da�x�NMT˴�����U�0��jl�������o���7XȈ&�Jh/�7ϣ��P���(7�F�_ؼ�pΑ42d�0g��vę�o�Ky��(�_fIc+\8�|�$̽J�s���mTP<�3ʹ7gW��Y_�#!����U(7��.Bv�i�����3�'oIX�d�����}RT{7�ӻ>,Z3f!�8��*�6���.�^l[�3m���O(jk/���E�"+���@�P�ra�)��~��������Ѵ�4zj2a���>!8�湆�F��L%/9��y�M����NɊq1SS�#�ͤc�ۢ�ZV��tuꙜ�ϟG�����@��
3�b���v�O��'HO��v���hWE�W�x���E�r}��$���t�Ǯ�&ġ��_���U�� ��ێ$`'T����XZ��+����硿��7Y�놓��G3q]�C�_iP�H�H�-N���r]����d���Lnj�!	ß_љ�Pt�g�Bc�ݶs=�������@ ˞% 6�s�4P@}�����[o�o�����,����q�A&��/���&�����z�6�=�+����	R4.m1����SЅ��U�~����9����V�L�>]8��u��-�K{����_U�n��*&�GrW?��/�����	fY��'�����4S��<��w��G�����u�OB�V8�d�]0����+w��3X&�(8XqԺL �i�n$ ���J�����N�a\����KS?���d ^���i~$N|�TZ��v	Up�oQ�7=��\�����ǋ,�&yu#P�?���jp�s���}KF?eX[=�=�y���,U��i8J���j2=�9W/�{@����Z=u�
��S�[�-o�{(z@K/���fh���=X�D?*Q;����4���]#m}�4'�K���?��ɪ�bR�g��"�r\z�s���w�|����0B:;c��tϟX��˪�){��mQ�Y��є�褕�R������v<'{|D��&��}x��Ii޺���%�w�&CYw����Mdm4��k�y�U[&k�9�G���H�hf1p=��%��)?�ߢ.�5g&Qp��K�0%�~'/�Q�J�4�_l2��j|�UG�#��&e��4[cA���Il��j���4�a���*�u�%�
#/��y�K�*��2�2�^����Y���Bf
E�-����x��b'z�Y=C�V�W�2��D�\ؠ1n�7@�CF��.��:�����ⅆ�IؓR z4w����2�3?��vO5�X,���.�S7N/1� �C�خ��0�Bo��͌d��ܐ������/ �V��h[�/�X�����J`�1B���<�O�iir���F�����z��J}dCV�=�zJݍW�nT��m^e��BH��M��)!��^
�:*�!�6��{)J��N�g��$37�;bJ�3��#O1ߵ���JR��G���3�-2kv�/m����\]M�~��IP[���MM�p��qd�3T	��s��MOI��=�ͥ����w>�v2LT4��"�ۛ(�5��3��m�˅�s����5%nu�2yJ!��ðe�z��>����e�׎����t`0O�݃uJQ��W��=�6�g.�_c4muvmS�7��M���C�I܀�"�	2��eK��[���0��Q鞀l,��lD��r��������E�	(9�D�,j~��d��&�3d?k����1%��˂������P]�
���e|�%�웫|,�B��1��@�c�2{ɤ����T����W>}�vrK��I��L��I��Q>�OfP��֖�PK�T�yQW��2o�	\���� 5�h�#�C�%�B5�X��B���,-ɵe˚�gB�ehg|^�J�uo2����7)�-z��5.���kMFb���s�c�B������E9��J�K*3��Mڹ/eJ�A���H�Ev��^��>�k4��_m3,8YZ��T6����{�X�j���S�^n�RmMO�Z�>�$PhN��,'=0�q������;.y8���0�r�_|�F���w�Ow���z�!�K�5������&Cft����G�M̌��M��8�rR��q28����i���k��XONU���L!ÚR��Qg��������j�S�w�S?���}���e5��6B�D�5��X��+'������ѳOd���4����H��k�L䴠=c3�N�W1�����{8��10ĿĠF
ʎ�
�݂3f\BL��qUK���v�/�8��)���ʃ�D�v��\"��z(���'va��o��?[���U��yX�DG쐡��?��'����e���g_�&$nGp�������ʬY���z��h9YmzM��[�{���4S� $�� ����HhX�a��zu���k��n���ə���ð��P8	�&��^�?98[��[|�2��ӽ�Lc]��3Y�>�x���`�z����G���Y�i�������d8��^���h�R�݋q^��Ѱ�HBG�7�,�O9�`|R;�
�?K��k��mZ�_XHM��e���M�C���OZ����J�f@8	q�A	N�1�1v�_s��j}�Z�\@�l;8�A`B�x<��`���'E��F���kNQ��M�UaK�����B������M�!XFsw�ń6�J��(���"�o:��<�P�"��)n�*[�D��W�RN�e��7#�j�3�P[q?�s9�A���ug�y'Έź��#h؆�ږ*�S�ō����ϧ1�-��b�����\�Oc��ߔ���\�*����M��_(�� �A0��ײ�$p	��;7��]')U*���W�9�MV�yA�Ը�����4�5](�7|4ߥ��M{�c=��˾��^�����=��P[O����:,
��*eAG/��{Jt�q@|ĕ�v��u��1�&���5��DT��s��t�j�Q��.�GB�JK�Wֻ(�^�m������D�qR�0v[��H��ԍ�vW<��h���N����u��b�EwiR?'Bm�����I�z-��T+f)4
�~�[6aV���ć��2���(�g0�u��=+����������/��ʇ���e�I�� =���-����٬q����{H��g�١3����۷��6�=��E$��0����C�6�rv�=$�q׭e	�;�sD	WR��9F�a�z���ɧz3\�|=�M�ɛQ��ۿM�S�iۿ�K���Z�r����]+�0ۛ`����lQ2%H�d��6v�<����t��y��رgԚ*�-Z91�vt�}��ң���dA��Qo7�������Lߟ��-b��+H؛���F"���_з��$nm$�Y��5��6|���f�؇Pc�L��>Bw��3"97���A�M�y�v��:�E��WM�2D��4�b]Æ��"
׭��N��$-A��R�eg��P��ӿ��2����a���y#}��:[hUǁ$?J;urcަ.����\�������c�� �_!�F2��:�?��6.n�Ư_���Oǁ5���:�wn��!�Le���w.��Y�4e��kM`mł�����c��as������`�Ν)?�Z��)k
��)7<m�4!b�>�j�2��s3��ʼ�o<���!ٹ�t�?��~НtXC�O���K�)u,K&}��$��\��w��]ءFrV�p\���R��!�b��)
I�8�k0�7�&��&������Gl����RBd�)ͱ�"b�TпQ�	1�V�>g��U���GW;/�j<IUM�����.�8���_���"xm/�9T&�3���ﴳL�nW���N�et��Ɠ��b�����"r4�l^niߵ�O��6����c���Fފd�R�܊B/��vp��"^��0��;aQ
��̭bװ��4T׎Qv�޴פ�X�}î((/�ד�\L47�{�ux8]�?h��$ʬ9i�~�z37��ӹ�f�k����d�� Z�2���/�j�^lp��0�1O�TR��eI���0���I�"�]�H�X�96�e{������X�"�Ʉ�X����T�x�N�~W
s7�e"�}���	30���k��>����_	A��*�1��6☲��߼_t����j#�L��=�mx4�̓
E���JX�͹-�E{�Xo����	�5��p���d��f�K(��9x�rYu&�߲�M��F#��[ĕ"���$�N��o��U��E~�����>�5s�%1Y+����zKT�l�~47u��/եy�.���pxw�F��0@��yk��&'�Ȉ�yzl�5��A�3�ε��+�ZG0݅�a
ʵ>�
���������˜�15�����Ϗ����@�*��E��%�1�è��#�!�p⌰Z��م�<��׍��~�5D���:L�¯2/�ׯ�QRg�(���o���ˋ[��2���[_� /�h?�"�q��6�Q�z�r��-���bF�NH� s��J�J�?z��i[�[s^�9	����+�<�!ֹW#|\6��ԝ���7���J�g{���~@ia;�?�jB��ˑ��8��]����������ي�P#�,wn����V�l*��n桾��������3;ܱ:6�#�w�(A���2<_aLT�`b��^̼�����~�TrǪ6P���w��V@��a�i�6m� 3�L���ë]x��D(a�'�-M���@}��_GDm���d�{#���UH����ĭ��a�>wL�h�:�Rn����7{u�zP^��ي^-Y�E�3EW����F���Dm��@v}fŶ�����;	O.�fii��گ��[�@˾�[S���e�n���/������{%?s)��V�W���y��ȐF ��%F��s�d��S�����'�fm�BYY�� ~̶�4j47{w���p�Il��-��)�!ܱ�h͘�tG1B���S&�O;A��rs1E�;l�&��c*������K �5�� W��.S��=�nk]�����y��?d6��zT�����x�PK1�������	�����,�m��f�u�W`�ѿ�>�S�uфt�ZZ�|-`�?��\s�5�>6��d0`
]���6|!��@'��TgΗ����Ha� �h��D�[��F�,~�ҜF����h��X��rX��l�+j�i�[�9���<�D[P��5.��MZ�v���`�>w�n|���c"nuAh|_3m<i|����.(�i*��cM������t�ţutK�~��p���c��f]t��9���ev0jL�_`�@`�f�d�п���de�nX�F5���a�H{:y�.ց���7��,[O�O�9��G��q�9���V�����qm��ܣ��f5Mx���Y����s9�oRk�y"A�/j��,�~n��F�8����M�k��bgI��w���>�~~k�G�H���i..�S��W�TvФ)�JcU|�R��<�o;�G���l>�K���Z��:�ŕ|���.�/��m����̝�UL���^��i ��n\��q��N!��{�3��&R̓T�ؑ7�&i�r��(P�<ƠP��]�4 �CƦh�2��H��k��Ki��I x)-��Z�ƌ,@g>������!�] �p���˘��)�
@��1�C�����e[�BH{iI�d�@SÅ��r�	��P��TI��4����z��z�&CY��[��H�W=s�_&���o�(����y��� �#���ᘳe-jUK�l���|g+�F����������m���>��G�)��KHh=�c�g�����[���D>���V�*O�XB�439���C�N }tEM��rV����a��k������n��I������guZ���r�����j�٭�J�?�;�J)��r��bi��L� ?݊(��ڪ>���K��[�*�Oٯ;�.3�m���F���Jshj�ڭ9:jt=����[�~�y��lĶ�����m�v�1�u	\�=�K�!�Ҁ�a2D.�g0zjW�xL��|�K�pO��:�褀��BZ3��^&t�@�ҸҦ3�k�[&������([��-��`���B$M�P�tK�zI1t;[��<�1�G=�Pv�vh�uE�� MJ�3ua�	���e{�X�Y��_I`F� ` �����wg�-4XgL���D�X w,h8-��q�7��?Ԛ�� _�o1�0�]�jXB�B���P�l�?�9c� �Q7�69�A}^�v�&�Dd�	�D�LS������r�e��r�\����#.o�&��w�s�GE,1���/����.���:V0��?Cv�y����8n/��{E�ǹS��������|�ki��;i�7��o޾3�a:��V�Kkŧ�gkH�iͭ�ǿ�y���쏄����f�&n�i^ QZ���lf���^'?�G״�2��ǗV�{�ּԂ��-�����;�Gs�gio 3'xl.A������x��oF�s��2���\�>̺����Ca��F��0[I�tE��4]BL�eh��8��"-
�y��~e�Hә��=5����{���h�hS��SL���e���PX~�;2� Z��d*����}H�t�a����^mkw������ޤ;���֊�����^`�������y�%�Z@���{���-n,2cq��q{<��/����L&��t*��#�c�o�ؒ;3����>;��U��]_�\֟>)iF��evc#2��̑�_�I..��@�)оC4���qS�2�7�����W���s�`�3
��9�3 2
s�	����e.�}k�6���VJ�u̝�8ۘU��J�f�h�֓-��������l�-S'�첯����=F�_�X1l;
 � ڵ�c�-0��L��{M�/��e��(*
�H6���.~"푠�5���?Z7�A,�����9NO��\[�|�H�k����m��~��׼�hX��~h{����q���%�V�Yj���ĺ 𵱶��Khm1m�M�U����K ���q'X��>���I]�U�V㌭�Ú�M���m���/���s2R�?gG$*[ա
|w��3�@�3Z��T��P�{��?����ᕘ�o��OK9 NL"F	�1�vy�2gۄc���}���JA���;�t�4�������}oL�ƥݫ}��Z�5��'0��(� b�Y�!��kLQ�ML̠��ɗ_�S�hM��K���-�8�<�gEf���B��:8P��鄧:���Ҫ�˦��1�Z2��4�Z�}�@����&�N5�M9�7Q��Q��U�3*ND܃���E��WzTУӱ��P�d[Q��'��s�G���E�/����� �w��Hg�NbK^��k�qv6�Kh����4*	��
��i1�����~/u��M�Wݡ��݂�-d�Q�V��X��O���2�x)�����;���@nޙ�Ĉ`�
�ڥ�e�5�03�v����g��I;��!����iF1@�h�.PS��';F��&�i�����+�ȟ��~#����a�6ףafN�DAz}.8�,Z�K��e�׵��'_�u@͈C�\3~��Jy0�X:�(�S=ш�>U�7���ix#M��B�̤'鳱�j靎��`_o�=��|�K5? L<:�S3xd�����)�k ��fX>X�_��>{s���������.|��I�Ϊ����e�Gf�\_��X2����'kQ�� ShR_�����R��&�J6����yq��{��]h�jQ��>e5���v�6\[X�*u�v`���γd>��t��^ɱ��9�@��(���#�G�v?�+:��c]���B[�cv��믇���6( �^�s�H��1�W�u�N[aF5��T�a��)�anu:�4��f��1�W���w0���G�Cࠍ$�A�s�8�-照�Բ0��_7M=�M,��ۘ���\��?��nBc���&6��S�q�r ��U@l�����ˑ�&a��;���"��T:@N�X�@'��,��D��^L�bXjܵ�!C�2'X�­�)�L����5��)�~���5%,x�*a3旒�{� 5���$+���K�x-�d�m&^�ɜ�,���ސ�� E� �3!h�zZ۽��q���{g��G�PI5/�����V���ky�,�+��\�l�=:�����	"�S���a6ܨ4���;1���U1�h�hO�7&F�Y�5�� &�D=�O�1�z��F�w�钠�$'�i������1��� ;��P 3u�0`]��x.LD{|���&��7Z<���bل�2�[+*�s.�Y���O-@��[�nROU�cx��}��@'Z6WL��kM���dX�/�p)_q3�&�_C�Ο��=r�L�4�iЙM��Tǜ���(o_k���nm=9�g'���o{��^� vi�5�U����Y.�ϚW�]��OΒ?�Î��6i-`�t��n�G�Z8����է�����k�ݱDl4��_k!���~f��r!ˍf y��BĘ��V���kK��U�]Q�on+�J���S�/��/񏛠�2������00�GCØ��%=*�֓��p�s��L�x�R�p�bT���P���O���W�B��r^i�0/����|��.}���$\ 8`�&��L_�C�C��2�յ���^5��
�C�-�5'3Q�D��h�=�x:��56?����j�>:V[&�k�qڬ.��s�8K��fW��m-�T�"3�zQ�"Qϛ�#'���&d��\����R� c.{}�3�SRv��a�
��Bgs;����Q�\���oZ���v���&�h�fy�}i��yZ:��w�)'�sXG�"�F�=	c֏r��vX!l5�w���vV93�m>���n[�_�:ˑL�1���pW4̶�@��;k�?��R���v�����s)-wA���u^������� �0��}D�� ��l�Dc�>iQ!< �p��]^sb�eB�*%H���( �R6��K��oy�6�)J�w
�4��x�0X��Q�AG��oq`�k��}���k3���'�=8��*�3jZߵxƔ[�΄.��c���@x�ֲ:8��	(�뚯QO��<Ƃ=�֧���-Q�h��FY��x�m�!ˈ9>���`qǷ��b�);�^{k+ _:6 �
kʶ
m�1�{=&c���v���@&�U~�h))늵YK���~T�����j�M&]�8�c�N%83���h��J(ص/��@��5�/��Ğ���\����~���G��(z�kA+�uSU�?Ξ��~���%P�C���Ó�OU�T�������"]-���1��[�\�n�_L�0�K�i�iP�.�i�mj�O��YV)?��OXڞ*���1��mW���M��V5#��[�4���:6��Q�D*�?s�����P�9e�3����B�*p����2ʥ�
�u8f��2p��/7B������|�?�lEw�~m�&�d#�e�H6�4z��9���N�L`�NV���Z�V��h0���c�h�	�����d���uZ������n�������C��#�}���L���ڷ=��H��s�	P�/.�Yi�.C˰������h9hQE��.X�:�6�B5�f��oe"�LW��>'
t@?���̅_��ZJ5UQiSr�W��n�yiր��[�L�tc@�;m܏�]k�W�1~��4S�#�V��g��:P�t77"��������+�����L�0�0T�-��8

������ 2a�sv��1rN@�S}\�Ń�0��߇u�Ơ�q�k�����\�zh�T [�њ�G�񚕆�`8���WB���1�f���Ą��k�����ϧsnB�z���d�q/�F@�{���Z+wR�����54��2��,v���X(R/�k֗�VIp�i��f?����֑䣖��#{�T)��kܕbȆs�
6�:��ھ.늾���A�怜V-����X[]�;o�k���\��&�i���s�@�s]ٟ8/��R�`�0����p{��Vb6����)F��<Y���]��g�fҊl����r�����[Ɇ�\}��L�P�m����!6�:��/�KQ,�C��K��W����6�������)�� -��hqh�~�U�`@�wԽ�Ý�AMS5d��Uj���S/�u�p��D@��Y��6?i4�0i�7�]�ܢQ��S4E��BO���Щ��y���π>��`N�b���-�C]X�~��WAWCrj��87�װF9�dȸ�`V`����)Z�m\-��WyV*�����5N50�8��7^�6ޢߙKu�C�@jf�g�A �'[&s��6(��`O�v�����9:�O��)7�y�$�)]�o�8	�ӎZ�{%�SZ	6z�A��u<G�ka[���ֶR��A�a���̤�<S
t@?Ӆ��Ӓ9\¼���f�Y���	�����\샢�Ô�VMp:i���Z�~X�J]t��b<��kx�a%<#��ģ!̧9FmPd�r��5;�Ϟ���\(���}e=X�qǬ��G0�� 0��M�5��^��@KU5ƞ�p9��3�hE�ᝯ��
����1�#꺝[q\�� ����hM�X���w�����ۂ)P8À�sl�j3-7@�)؊ :y�����/���چN,R"�3�X ����,�6cÐ����9p���b)�K�@�� �~h�����[Z����s��)(P��hQ�:�攱�@�������m\����%��^Ƞ��/����2�[Ӑvn�Ύ�s@f�8���꼝���䮵�*�r.Lq^�E
}�\���"�i��'�)	�B�k���������E��]۟63�@I�4�����)/��k�N����(�@@3w�[��0>c�0a@�QS�9��>����ۏ�[17WPsU1L�i��S~�++&m�4��꿠n�p�Yis��k|IGj���Uk>a�G����i>��Ր!p�X0�@� ��T}=����G�{��^q��'�ph5�A�l5�s4�2o��G�ܶ�ov�$Ǟ�9sO��7�	���scnO��8%/�W«��7k��υx��u����L�Z��s�-K�d��}gh�P�g�>ict�\��k�-~V�4�K��E���}�T1����_Ϙ��z�f�=kY��jO��9gB��5���GECB�|2G
f���YS��Y/D��J�J��W�J�L^_]+ڝ��ƿab�&���~�� aR'v�1T@��5�h�L�����~ /$6X�6c�1��`kE�0��8)�2���ڡǛ�eL̶�{R�昢��V��$�}9?�bL�O��cR \��c<M�T�ƴ�f!��Qpc�c`U�ͩ���5�x��	��v��]���W�k@�b�[`e��~�8S@�� ��%�Mg�����|�!Zr�Ҡ��DG�Ҳ�G��
cc��W,*22��Y\��X����2��qK@��D�0'�>�l#�Y�r��V W�����ڎ�
��X�N�P�9�u\KVH�e��-��?�È�$b�0�De1Mj9�k�=Rlg�^���5���Gv@��.ݟv�b&+�iw�0{�f��z�SX���ͤN��������V����_::G4�0H̴�i�Z>��GM�9��03߆I��
�Fӣ:�R�c� &a��䎾"L��ͥQ��� ��R#Hx�	d�A4��U3�ƴ��2��}��;���0f�+��㽯��b0�t�&4M���DS,p/`oڴ�m���.����YU�u�ZS���z-r�Z46=C�l�ܫQ��V��\"�$=�^��Mh�v���{E�̸G�/X3-�V��)M�eN���0�=hGJ2��;���4k���~X`������;i�A[�r���qy[�O&>Ror�K��gqC��߲�[�zD�~=Yx�gԽ��+�,j9Yƒ�m-��s�@�s\�?bN�?!nl#&t+_�L��?�F#uʍB��[�_�.N~r��(w󘴵'$�YR�:;�C���x>.��|�>"���E23SkL�@ΑĔ{��q����34s�kv�xF�l-��q �w4}�:R�^^�_,��%�l�$"l��8r�����n?�a�(��5�-���>�πS�`��%������m��6_~~@H_&��'f��^PO����Qƙ�|���nu�H�Z����\���+�jV�E����ɟ���g�Էm恶-AY�+�:Xt��%���,3�&09�,��2���*�0f�Pv���8��k��5�\;�?i�>�^������uR�Bd$��ZH�_I�Q�C�wWH�
�G43&�v�ϐ��pQ��){��޳�/��~�����o�;�ݗ
ޡ����1�aP��y�����2J�pSs��J�^7f��&�dN5�I���,������?�Q�Ol��k&�*����h�|����
`���<��Q���
kLz��T��F
 ��ӼC��7=&w�)�T!]V�&��B[.�
U�`c4��)F��o$\Q��ǰ�8g[�=���7G�#�ۯ��AKG����U�"(��e/_���k��%!�/�8t�e$`]��y�=�r�n��Q�w�2� V���h�l����gv���X��2�K]g�9DP��$"��}?8�$�ܜ������ǻ��IJ�5f�%��4^�б��j$���PB���̳d�{f�ښ�z� �4:V<�����ˁ��3%��<���f����jK���/:���������[��=�~�ٰ�y� ��Ϟ�j�հx�~d�6Z[Ѩ:ҥ�4�wmj^���YN
S3��	�W���2�y����)&3FK�%ÌY_�K]]��.D۷�5��`�{p]� �� ��WO�`i� �AOSk]t�����K���j�g��L�b��N�o���ai̺�s`
�/A��5W�GZ^{3ó���,j�#��"@@����#�N��"�D�h�$�U�������]�c�$m	���-L� ���i^�?���;7�oelk�&_���~@�)���*������+��b�J|�s���q��`�钆 �m�}"��ʄ�Ɨ5K��Ci��� �8=��$�x{���=�G�&��??��χr[bI�]�A�����ׇ}��k=��وi�`K���$c��2�^�p�ו�W�/���y���7������J�ES(���͜�0S��e:M��9x�aA�0�&$��i��U~f3G@�f����fЭ|����^�њ���E�Y� b�N,���e�6����YFKC�8Jϵ���HI2��=e}�����M�5�h���[���b��NM�'3|s䧅)�'�,�����-0� M�3�A��S
k��8 �����y�(�n��Q�7� �<��<�yA=B��!l�H�C��T��񫷽8;���w�M�GY$������~쉿�0��b#�M謅:�T�^��֝�V�l��~g���j<c�Y~����R� ��n?�1f�u�ߜ��.t�N����D!J����G6D���SK���9D?��@��?�U�w0F1�5�q�������Bu�)���M�tz�f��X�`�t�q�� �� @kF��`�ֲa��K�����`Q�+S�&9���7��2��UL����w��Lǘ��[��)0/fNc�ҀZ�R�%BJ�i� ����p��)�����O=�z�G��2�2��	�I��E.�]�̀�s�/wG$�qWDh�^� mt�1Hδ�h���Ǐ�F����>��BY�7@����3� ˠ���+�j��Ly�V�F{'�T/�2I����	M�pj��vQ��G��E�Hu�m�U;`=ۋ�������0��l����_Sa0B��Y��N�~��wpX���z�v�Y�N����.��Ӿt�5@�(�9�i��v�tJ���:=l�������� 0c��@��˩�@�9:���������������W����ޫ�ꓧ���$̄�(Za3���D`vh��a������R6?7?(�7��] ���˝R^t8�0e�uu��1�sUdt��wO^�v�Om^5?-�m9�9���`��ʴ����Q,�yE��h7��d�9��ct�i�I��q�fv�$a�BJ��%f��֔�G݋����j�-3��j������ڙ %�B�#(�\p�U�Ϩ��(�iӚn��SpO!�,}�1۷����q\�=ũ%�{���"BKK�K�CL��6+ݬ!x����[�(�up��������ww�^ ��H݉��S�߾�4Ni�ѼW�,��w!c�pBj�n�*�k�oB�!ƶ����:�l���z���}X(�DeB�?�w�o`W�����+�/�y�_j�=m����q�Ϋ�'��xX�ŐT-nؾW+�;�B�# nv|b-�X�9�8������l�ta*T��kx�Rzfd1f���aCR#Ә;m�ǵ���/h�ŀ';�8�\��	��y��&Z���GF�D�9�A��FK�5+*`^�f&ܓ`���� ���;wżj����{�x�e�,M�izW|�h|w�n�3��Dhe3i3S�Z�be.F2��F����l��[ U<�\��o1}�g�ˌ"����\�jmsjģ�:���9�g ��U'��l��cnw��B�hbp������, @5=%4d9��>�Fƨ�_3�֔Ә�
����Ecv6�[�iZ����lw{3�YTte�h'y�9@���k��Z�F�gc���q��0k=�<m�K�i�#�8�9N,=��~?�Sp�e�AK>n���
I'�.˗�!�t�����a��=.W�jC�?gL��g��?vj�����w��_\- ���V^���~���!.U��u/�q!���usV��;���ViU1��4��#c`�⏄��Hm�D3(�0�\�;G��KeA0P�v�75sy�B�N� �)@ &�C��s�ҩ(V�57���� -:e�9bb1�ܗv��ֺ�A�n������K�Q���í@Os]�X8��`=g@����%��8c��f+%t�K�륀�D�����:w�yތP�[��xļ�Ѝ�q6	z�
�o����e-�g�DnK�AH=7��v�y7���,�s��5�Z�e��7�� _�wϭ����m�T-�f<��l�F\-���pwT�$:;>k��������d�h�v�B�����X����6��s�O@𲏚�C�!��^����%��4GS'�B���M�����Β���e�S ��d?�}�%F{m6���KO�6�҅֬��/�O� Om~˴�A�������;�vM4={ֱ'�z����0kw�\])xC�f|�XF���~��w��۫�e����u@�/ޟj�����������L�� ����ڃ4
�\PX�Y⏟�)8 ����F[�4<1a�?�d?�܋Y�>��'�I |���ٷ�Y3�cJ�K���ɑRE�:Z�q-f8�phnGA-k�!(���D��Z 3� �-_s��P�E��l&n�՚�5l��%5���
s�og
�?^ ���<L��������-hRϢI�t��Rt��B��߹�>I4Zj��X ��֬��V�?�X>�|�A̷1Y;�������0��Wk����*�0�	�i�r~�O@���5-7 ���gӷ�cOid����"t�..�B��f���#����N�#�f2xm��Q�:%N!�}�v�(ͼi����̽���Q�bw+!L-u�k�|���H�No�^ZP\r�㞱�3Me��g!�`+� Y��R��v=h_nD=����Ŏ.���!pXv�z���ė$�M<q)��~s{�x/�؅rKx��f7P�O�/�u��R��?޵�w:2���Z4�|��	��AL�hF?tx?�
��r@�ͺ@!�#��"��VZޛ����f�."�G��QZ��L`�8�*�'Z�/���8��_K>n������d�u�U�&a���>�y��-�L̥�T�u�e��� v�j�W,�>��d0v�ǚ�f���wy/�ܣ
 lඌ��9�,�ɉ�Z�6�#$��G�q�`1����u��Fc!0N�ɬ?��R>z-����t�K=��m�W%�^:�IH)�)3u{�)5hz�/ Ľ}�F����{�1&{R���p�6���D�[�a�-�q�_d�� -�{�@�"�:k�c��3K�Վ�:��G��\�b�FL��W�L:��^c���t�6`����5P�!�𑛽�V�%���Ѣ�'o��A�]��#L���UA�>�b����*�����n.�Us�B��K�e�^���Ά����=���˅�M%,{�v���X�k[�c\�rϚ�@V�w�8���)�����NO�a�n6�Z��nmp�Z�8[�d������FdD6�c���a��_��K�(L_�a��=ȯ���M�r��H����~�������hA*��4�b�M{u����)G�iAb���7F��/2����FO��~ �w2���4'�������O:���I�kʛ�� ��zi����1��lv\u��Ë˟n=�g�+s-����D"�({b�\��l_���EW���w20]K���+]��ز��'@xOxa�P�;`'����~r���1K���CC�la���*���yXR�T�A�|���Y��3�}\��>�5�<�е7w�����a���w��H�jnvM�ۆ��]�e^`� L�k��-��Yz�K�����Tb�.�|!�#�����X{���fV��dY(Gx��d�W�򣊰��2��'P�Z�+����e�?��:����O9tG(���w7�Wnod�|7���4*Ƌy�!8�#&�H�@����H�A៘n���`�E�ұf����W�������*�=��.;i�����]�m��1��ޮ�U��F��4$#Y�N�L��F���{�&�V���-x)����=����Fs�����И��?������:�P���u�>����ǜv������X#����O���a����o�}�����ŀ�= ��R�m}ֿDf���<���"��W`���'�{��%nq�X �����m��\�-�V<����;�|�xQ[�5h1/*�	��,?塇Nh�qy�6�sh�e�ɖ/a�}�C��RH�t測7r�~�捾����iQ=ɑ���'�JK]�\�j��AУmB6m�2���z��%&�)�r�T���`�y?1'���M���O�VA�Z�G���lڸLR��Ѹ.D3�[�qbf���v<0V5f�?h=�!�����#:�����9}��߭������b����1��b4�bV+�9���!��v.���@81�4�$X��������Cl���\Rk}K`���SX���&���ۄZ&�E<����h5T �o�Xd�����Nz �x���*u�x�5��j�ٺ�)�e��������uO���[��eyأQ��-��?X���kn���ϯ@���]*2z��A�V{��@2��
��Eȷ%*[Z�V�yP�Z�`�d=0��j,�W'�/�K�Yը�-
��ҙ�����lT��T��Kp�}%0����4t�XczGsD�vʔ���S�(:CC��q�(��8��5D�k����'Z�����ͥ_k]T�֋M�d(��O��/�E�=��}���_HL�5>�(���;\C��B�f������+@]����a�s)����P0 ����Khe�
 ��5��j�eb_k�	w.3�{���ds���o�� �\���GR�����1,,D��.��.�SD�&)�D���yQ���k����vy{���7��K1y�3ϥ���>�_1f̺�@cq�OT�(.b �����h� ݿy;�~��p���#O�i|�b�bv��2Ko�GG�q��J�I�W���g��Rˇ��e������5&���s�N��&L�<*f�lb�6g�md�XN�g��h�$Z0.G������w���S�����@������po�JhL�@7S-8��u����Nv[EJ�����W�p����5�-��v��nm��y�r��n�z�q=�������F��B�ݷo���K��^&a�� gtZ9��^���M�eaIK#��~l��`Ks�9�@-y��3����R#7ʨ���(Zl�lh�e�9�G��'"�Ŵ��D��E#�1G�+� ��|�@F��cF0�8�r���N�)�4G��^6]��#KP�Ӏ.���S�#�Ki�k=�F��^���wI�$�Q������{�D�2�bbZ5����
�Z�]�F����YuE,`7���r����L���[a#���(���"��c�����?�>��j5{�~��?x����U�#`f��>{1����|ykK���_cZ�1�:�9��E]Єa򤲉�b�~+?��_+Ղ_^�G'�J�Y`>�6�A>�-fI|�����9�����P�WfD�����Z=�i��k�O�m�ֻ>��jvw�s[!a� �0H	� "C��a��*RI���|HQ�]���rHaH���a	c,�'�vc���"F���{��ݮ5�����|��s�Ͻ��{����g�5���?�|�O7�A2�Ȕ���%C{�k��U��,"B��9Sh�8ׄ,��Q��֏9L�G�b��V��9TV��ݻ���w�W��f�o�5��i��N^ އ�B��5�5{�7$�k���f	�}t����X}���0ٌ����D|3�ΧXHTqs\�;�ˡ�$��_w�	Anả�l݅��%u�����*�x馳�[�ˢ����0�I�֙�a�ωŊ�R���ѣ3�QD:;Q���<W������<5x ���,�J�k���d�ط�˺l�g���%�$sJe�I�cKˤ1F��xz�s��+0�vg4��/p~��CY��C��.�U�AM�ڧ0��֜�=Ҟ"tvF9c<N��^��\�10kJ�����c��n�������^e�#�Ӳ[�R����F��;��g�~����g��Z�/��d�;2�ͭ��;"^��bMnY�dRc%9!�t7H��X`�M�$Z>W�6�c��~حNϺٝ��-NF�,���{�T��p��v��M��T�U�4!+$B�Nd�=8w�Y��xq�Τ$��d��9�J�Z�ܱLE��B�m�i��d$�����&�2����D��Ǌ3�������E�$_��>�s��� ��{pC1H+���}��HY�z��*Bs"�>=��L\��Dގ;J�τ��^ʄ���\�dy�X���;/�s8éf:>�5�S��O��ͱ��80>xO D/�b��K^�u@?q�uz2L�mۡlN�>k�O�d��'&t�j�3�թ��;V�ݹ�~��P�/�ƞwd;,@hR$f���X�W�Y7��Px�h��Y/~��N�R>����'�k�S�|��P�b-=%\#�=,�
�14D�סk���%#,�S��9]!f�vނ��#�
���R����1!n��%�x��g�'"�l
��P�r�Ɯ�::]w��;���5��!P�~�F�)�y�g��t�����ӏ?�-/ﾲ���R����Ef���Aa�M6�9�crQ�U_S��;�M��^�u��t���E��G�Z$���r�P	��
���\e�%�a�eT[�C<�%@]\��T����s� C�;z ���e����L�T�ӌi�/^�dCR�]���n��9p��4k�A"&,���<�N�w�5�c��W"$h��\[H�D�|J���H����s'FLj$WQ�DʃעS�F�h�<,�I{Q��i|nP[��P"]����%��Vj�Lq�m�ý/|�X<^aQ�R�q���ٙH�e��Ǣ&���BAp�ObZ��55�Ei�|@�k�c{ �t(-���X9��Oe�;L�q���x./��l&V�ݺ���^�$�y�>t��^�~����
nM*j���7��j�U|�|����m�o�hBd���]cAx��ݝ�-��n���{cy*������ �H~��'��j���*
џ�"��h�+eVb�M�������y�/p�D7�{䇎�+nE�O�����"��2��؏�zs>],�������`Iۓ�<�*t�f������}�P6cx�(R�Ĥ��n�I������ !��e����h�i�R�r]Ox:y�����Zn5�m�#A1����X�d"� ��eMtΩ���c�R�	�t���K2�ǘ�S�ߢ�������:��%.�W����������e�@�'k�
�X
�K�!��*b��Y��l$řЭ��ԕ���A�HQ:��̔<�G7t��B���՘�r�5dzYd�]d`g2�Q��#�΢��4�,�-��t�*�ae���AJA$���ۚ5gQ�%!< (6x f�|�;��x�6r&�O�w%�QY&2�!�V1	i�.P���G�؉˳��M�1nV^�B��(k�����~��}�3����1G\��)�YQ�L�<�֍�=��'j?��.zB-��.�GBw��M��;��7���W��ǋ�}(v�	��z� W�J	ּF!�.y(*f����ѿS+õ�9��B�{n(Bn��k�|�>��MΦ���="c:��"r�,��)&K���5�;�m�d��V�����3�^riN"�����%�H���f�nYC��VW�^!��z�Ģ~ma� �R�Ѯvk��{m���I&� ��t�#V�_����1�?�*,F�	��so���{b� `@���Ёn!+}���b+�.n/�X�GVw�q�V��r��]���2V�#%p{a�0XAFZ�L	�8�k��l�3�e�N�sZ����"\�$�a�V�&

��	��g��7���bx���Bn���F[��q�5��;֋�����Q����t�X�]c��Sc��X����?�$����}M/��E4�Pj�H־$�+r><ޙl�B0�8�%���iQ�=	RW�#�b�w���y3��_���}�U"0�؁Τ����51vx�3��{^2�cM�'&�(���RFHM�k^!�{������#P�~�x����d!ޱ�I�������#�)�  �PIDATX3^>���)\��͢A<� H�V�I@B��#D>�0�Zm���Ƃ��5,=��aJh')%�#Q*�y��
��$	�Z��#�|��������?���
c!�!9�R��j�i�TC��~�ʀI0f#������"���풳����Ѹ��B���Ê��m��ÒG(A�a�a+�k��״5�p+4�H�m��#�	�އ�R�C�&z[za��q`(�a����������Xe��cA���㈥io	����msB�o�}Y��0�m.y܌Kt2��s����5c��+>3��y���n�>���*p��rw)W���T8g�>�ts�xKh�����Z)��x��$�A�a���^t?�"�2�_R�T�7�ħ���d��>y]P�~G��*���'��U�5�c]�x;�Euc�e1i@D),�S�إ�@G��	�7��B{��'Id����3"�l��ױIEX8Al��ƩY¸�!� �$�$� 䌁C�@���[��a��yd8ӻ �pO��tQVR��{�m�FX����I��*o���>���m� m&6J�H��ڭoBL�23�U������Xw�Qݭ�ޟ���.����(�'?.k�	�B��U�»1����YxlZ�Y���6n���ek�M�.Wʶ���#������{Ԉ�p�z�s��v��J�D1�E�4,�F�����1�˖��QӼf���3V���1��P�lm�#ӼD�yv,���W���`�g��|�M�J�*����G�_=�=E��~�:�tY��p6�qR
�ZvRN�[%;kF�c�0��l����܆X4w'��p��'ėm�B���\7�`�DI��mn��;� �#����<,��|��L��$bĽ��~���h�ȇ�g�h�{@d�Ok%O ����#X�%�]�K1i��dh�H2oK�����A�\��Ks�Z!�a���x�Q�\(S;o��-�K;�2J�V(V;˗�s�9���:H��k�a�؆6�C��z���K�\�|�~�;��.G|=��#�<�X$Q�q�]�G �Ք�о���y�
��xb�s^8KB�p�6���<x�aι�7��!�PP�x*g;��`�l��)�y+Þs��pux</b� "��7�m��b��FΊ}A�x(BFy�G��I�ժ��QC�E��WOWe#!)����4��B	a�DG+�j�c�F,6�־gӰX��vf1��K�K�36����
���n���!��xi����<G�6db$&!.�w�8�$ֳP�S���\�MGH�b�0�&�m��G#�3���3=I&��cj)�CɉvPJ��)��$ͻy���G�I��r44-CKu�,H���8��c��{�:��\���1�q45����e"��=g�"�����:J��d;5���b�b첛�����3VmX��}��=�����g̻���d�n[�Ϸ�J�%Ǡ�0�9V'8$[��Fh��;*v�$7F/�lL��QhJo��;;�=�;�����2w# BW��X՗��"��1���	Q% k3P�F�!�ck�~����"!���G�3.�2�ՍK3ʭҤ�� N��+�ĞLP�]�p��t̚�,�v�wF�$M��ǷAn�8��ݺ�8�V��7�������}��"j�]`};��J뙵����LQ�1�>�F8�)3�7$�q��;��_����Fk���$/��d(.>��BP���������pǹ;��1�7�>��@��m��}/��xo%+�r�t�WD&���zU*NV*�Y���cc�� ���Y�����T���b|���.��V���]��u���f��7�5j1�J2v��� �w~�.\��ҭI�Q �@�JR�����W�$���Z{ۜ�%��sމq��w0?汈]I	Ol^�~�(B��i���x��f,݉Ĩ\&7��Ħ�Ll��:�'S��K#>�吹��`X�����N2��G�/Y�E2���If��f�e!�B�Ͱn��%@$eq?����;}nK�����9���|o�>�iX��c2I����%��̙�-�/����ײ��z���-֓^S�Μ�X��N�s�������R.������K#w�[���u:>�W%�n�0���sa�o~H̬T�mX���F=��O�<�2��W����jI����Մ՜d��)WVނ4�O�Fd-���=��d.p|�� �;p�Bs{2b^�@PF��%t��Q�vP�������(W(1�q�8���|e��ʸ����S5��ع�9�R�h9�B�cS�h�L��(X��e�Y�^gޗ6�uM����G�����a��5K�s˙&8� A!yI��D�3��x��B9��B�!�Lq-^j�.s>��Bl%ʽY.F)U�SX�jj�����q8�c,�c9X$?E���OJr���H�D�\�MHsQ[9f�g��k�H"�*tW?(Jb�����6���Yl��@�a� ��܃c�w�2�˻;;e2�20�ef�g�#������|�^ �C*T�o�"�~ZސZF@bn��Z%��W�����Hv�`菓&�|�Wp�9��B1�6�8>I�$����Ę,&�����}ʎ��V#�$��[9~���Z*�k��3�3��R���
����7z������t��������<c�D�c�qG_�%����Na�3<f{�+��T���P�C���z�*j0ֆ��_j�w��n�_�}zzs�l!��$	�`�#��
�"��lxM����o
�O[|�:���{��٥J�Ui	K��t{%HY#acyo��, ,�kgd�GVv�=���6l�uV�M�3������?�M�wo��=2���X�"c�u�Q���8kO���ꔥ���V��Z�Pp����~�Q�L�ZWg
���/i�������͕��.��#�E52�0��X��$ץh��'V^�ϔk����h"ĭ�I�`;>�[EW���X�xeG�y�\��<���u�X�ޕVW�G٢��}?��)��%�GΓ?0fq�w��A)߅9Q�֩� ۭ� h�y��%�"c�|�D��ewl���y<��c�R���@�����뽋��m��������>�2��y��� ��E��nH��!����ҵ��k���4-Nd:�)��f ���z���%�ATǍ�a��L��YT��TlZ�B)���ڰ�І!��U�l�mF�b�:����ړ:)&D�W�d�[��f���m��8��N���gm��LD�������b�Gr_�o�Չ6#ql�o <�����ݲ'���(�FL���&3*�B�|\�{q�>U�II�v��I!��}S\x��`�:	�ϡhn��������@�ɣ���B;�r��e�Gm�凱�w�O���,��iQإ7S�<-��nWp'���Ғ�y���ΧT1Zij�T�<�uK(���ºǰ���>���J5���	������P��<��m�k�N��1�9�҉2������n��U�D����@�P�!c�Y7�b�f=�=E��~��;(aHB\K)��V���1���1�b��&Ă�ͫ�S1����$����%0פ��+d�$�ڔ䦶n��������,fl��]�"^/��k逎6R��)����`���|�D������26)
�u�{�z FY?�*/�N�`�:�X�d�� H��\�L��6�(����埪v;��-��&5�Q��Q"tg����x�L����6��]��s�Uai�n���LkI�V䚆��[\��ۄ����!�1�.jd������r�����O��)�� {��8��d�p���9�O�Yi򦥞�Ůu�-�hx�ra��4*�]��
[��6z%�߲'��2nR��ڨ�X�B�]��/���c�L���!��h0�	��<PD�~���ὲ�7����-'T�]�� �QǺ2a�6P-y��~��u8����@��=~���D;�mܦ�,m!d���Y"�֬�㭹=q�^��'�59Ć,v�<WA�R/�:�K	QY�ė��.ϴ�֫�w�7�4In�M醝�TjS���Mf%[�)̩����"t��!�ӭ�\�q�Ŧ}l��$4Eb_�"Q��/�*����XT��Xj"9=7z�Dx��ak-O��%�"��X��#�W�.�D�\��0҆��RО�<ۙ*���t+T�
E�e��%a����uÞ�b9�6_j�K*$�ѧ�ØV42�l�� �=���Er�c�,�~���r!�g��A7ۅ�&�bG��TcK��D�~�RR��0tA��*H�{e)�ҺGiw3�Õ��t6ֿ��*�� X�:0w>y�)�0ar�\�9�r�g7���W���L$��}Y� �e*%l�B4�8��c���R�Q����j�+F�]��d�Z}�~��qΊr�����O�:ފ��L*�1Q$�=�p鷻^/Ƴ��)*9���5F����9i�J�4�;�J���ƻ�JcI�i}֠��2���Y@!p��B��:�h!�� �I4�$��=��YK(.D �s�s�������-^~�n����c6�>t%/Ju�;����fd�Ǧ v
��!)��e<�S�G�p�}�n���!�o8ܖ0�GM'�� �ָ��Vz�Nt:{�yAħ����n��_��-����V��>YO��%W�����X���6�}����m5+\�"� 6��r�����D����n�W��n��bU �M�:����H�2D&tf��خu,bފ����.��+\��nNnk�ni��s�[$��&����n�࣮�Wef��h���}+2����tMB:(@x7�l��v<*j����\�����i��Ǣ��H�kq���"]J����9WAo7l�;����O�m&*�0���fg/ui����+�\�t��4n�٨�����=��24+��Q����Y�L���Ǫ
��[��|������/斿c�jh�mhx��PY'��D�='�BD��@�O�bP��v�Y���L޽h�-B�F\�5�Z��^��-(!�	Y"��e�M;�;V�pȬځ�5��>�mC6��c�.�U�eэU8�d7��\ �g����>�;�=]���C]�A�򆲍o���0��v!�b�z�V��i'wY���E���	"o�N�������YM�|�Y!xو�8+���IGWW�)泬k%�u�8�L$~��7����n���J������n&�'�q��7���W�?��n������#�>m-aK	`�5Mh<0�T,Z�Լ�^Ɩ�4���`� 3��M�j�0�P�V������r;O���u���~���7���;���K�)�bJf�Z�zԝ=��]����޻'^�֤�>u-���Gӛ���ehƭg"�I�#�Y_BH(iXܡ�y��!��c�J��{9�&M{��*N#7�
��'�Ǆ*j�i�x1 O�����-)/��/��46��˓[]w�F�Ѹ�h�-Ir���W�=�e�5�O�&���T��w�s�qȡab��S���~pf<���*Q��I�1�����_��}�s)�-�w��al�L.r�1��Y�W���D�0[�.��K��E�B�l�BElQ2�gպ �w��2�o��fw��/��_�6�/��}�,@=���Z�nm.���q����Cl�^����x��u�r����{|�D��[�zF��?�+H����X��}�'"�[i/����;/w��^��AJ��uk�i%R���ra�����|d.J����mouc��\;���k���=���g�6���8��{�&�Ĉ�U���G�om�����/
N�*�=��M��gD��r�o����n��	��_{�[���o�B�	E)W%0�n
����m��[�Ӗ�������g�Mmp;_�<(��K3f���k��u��X�I1S��QxS�s}`*�M	Nז;�j9���Hh�q(�������e.���l���8>T�����ݹ��NJ������X0�+e3<&��V���V�;ceB��xm��a}r`�e��IlO��?�P��P#<�??��u���:����2�x�	5��L����YE�h���	@i�#�l�ŗ]U΂����a�G����w������[�雯u'_�B����n������]�k���J�ӧ���U��2(v�&���5��X���N@1K�be�l�L~���v%�ES��f��H\r4��Vʸ�T&�J�7{Yd�y��|%�/o�K��Hݗ�ܖ�7��܅5J��+'ұN���c�N����)� Bg��S5�K�Ȝ�um�|�4��n��{�C?f�{��-\<'�#۫�u/2em����[���_�N��Ů�/Et+���{�&$���%����8w2�ܖb�H����i����R֏�q��2�K_�;1v^��@+��z�mr���'h8�Fa[�I�����]�%@��P(�[ǎ|,;T6��ų��a.mt�N7�s��(�����ugR<�"�ՃG������~��Jhzt�t�W��l_¶��Ieb�"�4c�P�����^��JOa�$��L
a���$���k����^�-Y�AM���2��0��Jvó<�n����.3��>�y��ť-Z3�K֑�犹n��^���v#Y}����ݍ/�%8���R�&���,ȴW��X8Q�Y�̓���]�i}���0��X�EOU��o�"����>���M�e�Cu�nb�-�@�We�;A�L�+��?'e�W?WR�U�])�jy�^7{t�۪(�B�v�Ja٪�[)/ʆ�Gb+���w�t��/w��?�����U�HR\\&X�j�����5�tZ�ͩnr�8���1O��	s\[��D<,+�n	����7>�M��{��+�u��/�����Rq��{�&�����\
��ѹp9U�A����>x�=| <u��
��=7njtP�j��Y��o^,uD=|Z��}�?��;��^��v�	�s��� ]�`�������BIr�W���՗����r�HQ����Kq�ЎS�����ǳ�T���
M3\�VV�d��lK���^G��AQGKxg�9s��V�J�~=�K�,Y�TP��j���1�D=�3��?�������J���M�*L�?0a��Ɍ� s�e�b� E�'҅�)k)����Rϕb�g��ڝ~��"����Rem��,p�e�����"�i&�P&�+m]u�M��"�|<��&$	s�h���,��2�́Y
�����Ӏb�hR�,4��Q6"�ѱ<sY��W�t+-;c��,ױ���uk���{Kqr%��Uɠ�L������~�;QV�H7�f*r�����<�(�c/�T��q���&�P��i[L=�:�����wS�1��@p��:�𵀏\�j�W8�[��z�Q�N�O9o������R��Wj������˻V4Fg
��2W��9���X��������K%�=|w�͕l6Y%��v}�u�d9i	J���<�ϠyQ��핯P*�*�B&���y�ď��$a&�ۉ�J��� $#rm�/���\<P��RDm׻�g��@�Zf��₂D8eL�<��kB+��ޅfu���vr�5�n�|���}���}񾕹K?<,j����R/�!Y��@�u������X��0��s�I�>�����+1��HA�@�D�W
$�:��rgJH.�]ߺ����L�c�4����l]ӎ�2�q�z��Dd>����@���+vtqmK��COPls��6����E�&��6X�c}�~���Ŷ�(7	Z�5�͵�O�,�ӗow�k��"�|{_�����׿ޭ�}���N7����IH��Ҷ�]Y�Z"5wіX��d%ސ��vw��;&�	xP*VG�XYq��1lsj�s�:k���P��j�PHx
"nLv>���. !��!Ғ���ݬ�,Q��䶹�@+�S����R��p^Y�ke�w7oK�yY�h֔	��On�t'خ">�Tcme>�r�7f�qe����$���_�&?�/,�f���?f����3 �!��ɝZ���.����Y�2���T1��kot�"t������ɢf)p3��$����҄rUcz�u������~p�ohygM=��	1D��R�q�/__>��?����[o�'�\�B�4!`A��u�%|�K�ĬLx3!4��1VAώH��ڒ-DUu."?��_Ս^~I��R����S����|6�Z���ďj�_]��!e�@�e�vxx��Jx���g`���X�Y^hٔ���O�w^K� ��m-�w��"N��VhBNu��f$��!�w��0�|�+_�fw?�n.��"�m��Q�2]?	(�+}��{�zn�fʍ�_��w���<T��{� �����B6?��G)Rc��fb��W�-e%����\�J
d���������/��M���;��2}x�q�$.&��(���}��r.����^+{|&�gõt��^ֶ՘` {e�󠀥ri�ŋí�x�M�z������g�H�K���9^�sO�y��'�j��Ș�2[��]`F���������_�f_�R�!۝M����i��e�E�RN�q����"���2H�����5w��N�j�Ǯ+O~�JmX�1iQv;:jg{~�~�@kx�F�q�5��?k#��n���ɵ�
&E��a� ��]�I��s	{�*�a9J4:��؝���X5��\q���˲�7r�.	߿��g���Grq^��ou7�*�-Y�v���5��&)��Mh�R-��JB�lm�E�LX~�A��eۓs���b1�&�����f�8�:��nM�o#�0׵�����hM�����{��� ��ޟc�:T��yc$���E
"xv��2�*>;��>��w#kr��T]��H'�����HQ�[B�
:�s�X�7��Z�ZɺV r?	|j;֝�Y��"/������&�������n�p�D	r�ՙpY)���s)�?�U��x���NS��Z��3%šH�g<�C^���"s3�!v1Ìv�gH�!>�Б��Bk�qvb�~�+��̘�a��t5�X��+"'��zSr>�y)%�}���r{���3���`ٚ�M.Gx����&vsm��ߏC*�9�BvT���S_~�u�N	Gv@��;(:��|E--�ǵG�������c���7lB[td,/�6���A�Ibu�f�_��fk=C�@�^*V��q=}>U|�KTEI ��K9`e՜�v�U��U��������ro�
��&���k�e���z�\��'�L&�rR�5�IpLo	J>'�:qZr��]�,J�T7I�˰�D�o��TT�H7U�$&BF�n�n�/ީ�V�b���zbm��Aގc�B_*0��O�z��D�wA�{^k����g%��^չ����Qƣ5����@��|��V���i�D�=�_i|FԐ�J���n��13)-��H�6�VK�T�ۈؖʕx��2�>����<K]�D1���ޭ��-��w���Dȭ��ZSN<[RJ�U1��t'�5%�)P\����_/U��=��
	�,�D�%�ױ�O?���Ӻ���J��[��t)�2"�C㶹��Nz7M�&Q�oJĚJG����<��	�|�k�����;�/�����]i���z{(B�����.I޹Pj�Kxb�d�}�	�CH1����%��X�EG��������0��:D��������R4E�؋>�*���b�c,v�D�d.�޼����g-�.m*Xb�2ۃ�bI
H� F�1Er2|��3Qa�G5��a�N��9.�B���o�ŏ5i� #Y�ˏ>RETY���Ն��uY�c�bKƢ$��6���v�pg�j�h"J��FY�a�U�-'�x/	T� �t�~G�Ꝝ�^�O�.����>yT�{�DL��L*1.Dպ,�����b�|�A��Ϻ}�O�l���W��@��\���ȁ��4́|!,��jfY�΅�pY�L����G�<�������0ѯY��|}����[����¤E�<��}n�X�>"�uE�[���{x��Mq&���j-���K���/t�W�� c@n	RJ���h���^P���1,_T8hŸp�+�C�W�ijS���i
����?���>��s�wѣ\3c��
@��[�Z��@�u�A�$H���Εp�V_�哛тW�Ȃw$��#R1$K���I"�u&]�*��Ͽ��Dű���k/D����G��=�׻���H&�����Dv��,q�S�U�u��dk�OD��H%j��l��5���k�7˚f�%�Gf�{o�4b�D�w}`$1�5��IMp�v:U��F
�J.��Zb���$�WY�*�n�+.\���V�2�]��5�!��8Q�|&׺]��ZHD��iE<l"�\�Ņ�,U�]�2'�:�1���є�Fz��1D��x��S:�����������)��tT����+�}v��E.˛$7��l�ߝȨpd�J�*�b�+�
݄��R���jv���cȼ#m�Ϙ����L�����������vͳ� %
�)*١X�3����{�D<�l�T�utGU���n�%U*�ue]�X���t�GW����V��RڼA���_�ށn���.�Pj}?+^Y��٢���,����Do2g��@#
N~� �I���4k���3�P!/ee��#P�~�Gxп�/R�����d�w ��MA�f[���Ēt*�$�$��Չ�E�8���HY�k��]�5VX8X��z���b�!>�e@��>�빬o���k���Ҧfu�{�c!T��y�5q��9�qh��x0e�}L��d_q�c�A@�ϗ��e�������n�*A������f�D�E�I�<Y�$��g�R�a��-��0�[h�p��\��!-$��m��o�����> ����]L�d�J�@���>��sa�E1В��H��QΔ���Ofݩ���T�'����$˭T,��� ��uw�2%2��������7֘��@�>	���DB\%r(�\�#4a�����e�P�2�'ZFy�/w�Wn�B�J���[���V�(\0���y�b�U.����v��T/�A�֩�����hRv���Ə��w?>{����m��J�3	��i�,D�L셊��A2z�:�#3�>�f�_�}Rw r=Y!�K��GFQ�^@��D�2�(�/ܺd�n1LpA��a�3��eNK
a�-f�&�N�Q�,DV:�g��X���R�j}Ｇ-f�át@�.:��C��B@{
oB/�����}��g�38.�FR��bi�7GI<���l���<U�����	�,)����+l��!�>�k���LO��R\֔�UU���?�`�{����� ��� �0Ƈ�܅���������<1٤�J��f�No�m+Y� r]�����Y����.SD�Z�8��\�ʃp$�B���&%=��ed�6����p\z���D?�
9WM�1�-��[�9N����7Թ���T���PG`{CIoRDN^���TK`LQ�*�=|����7�Rۖ
�k���{�����ظ]���G"�/`5����\��n�?A�~�*�'}��O�"C)�o&�%�>G&s퇾7��"��;�W��^�+1f����
/�j�czY�2'�i��!�m��`$G9c�����+��tܱv���-~R��-'�Z2����t؋:\��4��I]v����rs����PmS���Ӳ4�b�o��)$'vi7%���	�L�����&$�A����%�V�>��n3M����$x��/t�7_�:mUЃT�@V����*F�P%f�x�4%R���}V�v��>�
��|l��˽�G���S�ر���)� ���rew�YnA"�����Y��"�_V�A��f�9��\��X��,�i�T������F���t&��Ò�>�������>�VW;c�1�,�"�P}tN��n�����*��z׽|�Ir[�s��R=�_�z���>��B@��cp{��Kj�)\g�+=��җ�e�YٞB���b~F�bG��z�O��b#e|�^a˟a_o n��uL�z\{�Я��:�ZT����z�im������A�� 2ĲaG��+ޙ-����\��&�Ƞ&�j�դk�W8��-�����4�@����~�z�X{��e;��F.aC��f��G�C7�?��|��7�c�:!l��44�����Ho���Dk�����ul�c�� Qp8Ǜ�h��/˒U��vn(�{����� �Ǣ����;Y�OzP ������S�s?t���Ox��c�]��J��7��������o�"��\V��m-kD����p�}��y���aOx[=��fb��`���m���q��y��!�I`�;K�]����)����˯t�/~���c՟_+w`�x�]���W���9J��dz�d��"�5�{O,�?~V�,`/uw�ɕ���Ż�c��֗���ׄ�z�N|ɍ��HW<͈�X��1���iR��@��㾇s����0a���8t�:[��,���/�3� ���a�A������$Ql���zgfy,3��Ϛ輶]ސ��4�Eo�%���$ɇP�� ��kb��� 5�7or�$�C�q��:���U�������-��>�W�$�i9T��7���~��	.�I����*	�x�TV:�����c�y���_��$3��=���B����5�5d���}��O�`n
�̵M��_�w^3�+^}�j���4"$�
��şU�f��]U���E�J�w�Cɳ����c�X�Wno̕��7s@�&��59�qv��N�dK[��U�u��:��X��/�Ax����_�j7Վw�kT�R�3e��@�<�|���{;V�����@	u"%�.���n� w��n��~K��!���l�~�I*�Y�V4�B�ǋ�@��0ʭ���#�T�!�0�oFa�[�M� G҅l��O2��<�(�pv��q~k�-�����kQ+��/��-B���m-�~5S���X�vЎ�|L	p��{��l�I��>����m��I��F��߻��|Ը&)~��ؚ��Wr����?��WJ;Q����~�[�r[�kar�z�/��a�T��N�(�I�d��G�2�ɨM,��;|9��v��A�
a0�4�������D�9f����K[���2����ǲ<�ic!�,b�Z|�|(�#ؼąw_PU��&�9{pt
��#Kcqw��ֵ'4�
�����ؓ�9�0�"e�$+]�ꂤ5iES�
P]|�V+��o���PQ BDRƜG�7� V޴G:��D�_��5�����������v�k_��5M��3�w�|���Qοȸ��y��+����J�������"�k=���{��������_�JjT�7%ag�z�)��ά�X��;����}6ZW�L3@z����kH���i�of��5�y�S%���I1εܢ� ��9��Eb#-���e�����6TZ8��/v>��I�52/�}��8w��W�%G��� o,:����6�3mũ�b��r���Kݒ����TK�ƪ��y�-{O��C�k'��r�n�uTo3�����y* �u��6 G����!����|O��ث��BN�Rq�N�f��R�Kz�X3�p�긍\�k�6��]�v,����I�q9�	 �T�T�sa8��$jn�߮�@xc��8��@1�����Y�G���O_{��d�&��T�~��{�S��6�����ld9ba���?S���Z&�q�9K�6�a��ȝ�񞣙vi�[I2�ѿ����D{n��#�����Q�Ճf�3N�G�����LY�/��/BFy�G	���Q���e3�	ja���ŁHl;ֆI8�:�0dJ�&��bN׷��	'���Z�n{Z1��uʕK9Ԑ�d�S=MBTӈ�z�]��}XB��C���Xqy/+��{nz�en��B�	N;����~^䰦|*%\!���k���W���l��VF�%�,�K�>�P�b����d!B�Ч"��,A�!�-�%Ǌ��&c�C�=���!l�R8B���6��(�[�6U`��d����M�}�q_S�,o�ڈ��R`d��雯J�����)��X��N�*j����àk����w��]�1O� h��s���D>���^}�;ז��v%9o�һ�_׺��~�}�Nw�H����C��+���9�gw;����nw>ױ$r����ruE��.�~�rD�ǔ�?B�n�A�ѻuK�+BP�{�x:�[��^K�Я�^�)��x�e��ڜ��sr��n'{Z�v��m�7,�HW#/�u�/���|�d�a���L���H����{�v�����~����Ma]�J	nS!�h7�l��C��"�Ҵ%�°��cX��/�����rWO��1�b�A��X��J;\�=ۡ*�<������,��i�½�;�QgZ㼖e�V����"�*Ԣ#��P�k 
iS�~i/�
��Q���[�vn���W`��7��ŀ��6(̉(_�b�h.�� 5Yܫ�d�R���9��W��[���"��{�$+�T��B<WB��_��O�y�H�H��6�Ao�f��3a�6G<'�_N�h
f?#����C�W'XĔ���1Ky�#��s����,�η��K%�-���n�����W�z s���-��)��2��O���8����zɟ� �z����>��[�`��"z����ӯ��N@3p�sJ�=�?V�xRp&�o�dL��u�z\{�Я��:��W��d�+_�!"T�y�p�8�V5�H<����30���;,{��ɬvIo��Ȝ��6[.Mh�f���hǭi�5;���]��oAS�w*�!���O6|#�=뭉�F�͢x'��z��C�*�c%�Űab�^Y�ڀ�.Xؙ���vw������������{�@WN7�/2�&.������#5W֫��̊%P#�@lq���]C_�gr J�Fc�٬�C���<o��p?'N~lsCc��.+cJl۪j{����F�ך�M�9a��L�	��R۩.��>�z�W_�n}�9-?�ƻS.m�L��Lp�m��R	}jg�LMo�;PҢ�V��B��m�������2�_S��#��Vu����u|��t�`96�1�w�:�* � R��R�ve;NaY�xh���{�?�����	1VQ鎊���1�\r���`��آ�O+�nc*<n��KWȎM���yF��y�O������%{t~�a��1j!�$�\��i�����Ē�	(�z�ܿ��>��eY�/�]�����7E|8!c�eIq�#H�jU_�RW���N��r�,i�u*,湴�w-t7�k�{>�i�Px�n�Zbr�C(>���Le\�J.�٫�q�_�.^�&�Ԯg�Й�ԏdn�R���w��ع��$\��Ε����v-�@ˮj�䷣������.��F�5�V#Ia��F� ��F���ku�bc&���T�Q�X�;�^�}���_�.���
�l_c9��e������䩎���x��:_2�%�Ņg c9��$�;&a*9f���2���͞3\��ݶ��oT�f��ݩ�D�|Em�g*x3z�,t�, GDō�k�#nU�W���.'7��A�wr"���P�.����
��6��VќգH
��� !��9dه��1�9m��G�d�a���pL��{S�S�X��b?Ù�b�$>Mw~9��.V�E��mD��Y%Z�����N�?uF���7[k:`kn,�c�u�A�G��%�@E-Y-~�-�갾�8�K��ύIl�A�(��8��~�|��ްDB��9���l��<��\f6� ��k�$o��e#n����+��P��	��Dr�	T�r��ݺ���F�
\w� p@��F7��JwS|L?�EX9���x���T��S�?�(�}%�|���]'7�	nv�(U�[Q�ԛ�h�:Ex�޷z���ۊҙ ��qH��>4��_b�r�6h��J��e�4'�����*���U�����c�6(�]mu,[��X�~�}ѥ�-U��l���� �R��s�d8m��������ǆ��
۫j���
7�5�T"S9sS����+ȋ�j��^R(,�3B#k�[w���ں�5�a�?-��-��]�5t�֥/Υ�����nGN���Vb����n{z�a�1��	�S�O�xY&
5����ڪdMj�/�,�S�D���5��_J d��2^�i�3H�;�̶!�_?w���R��������	��!�v��|��O����"��2���~�ZPB��-E�ls)�Nd�ΖQ�B��ݷ��~gR����Sl:�Unj�����1���T��H��՜]�½�D=���K�A�ؑS�א̲�ٲh���A�FX0��FQw\C�2���Kz�)��nߞ�vsev�^�!73E>N�Z���8�;�L�[��ܼڙ�����"V2B��P�+�	V�e�>�x��o��d��=����`��h�����Õy��D�2É��X�Ĕ��u�em$�"��ã�-gB-[�-��}y#D��R�k,d?��%%R��[�H����3M�%��_�y�A�>&�7�GC�&8x�u�TFJ��Eħ_�z�7�f��6�%�aN�T�]�^O�(�k��H�s/̷r�_*�a���^Wi^����rNh᦬v%�-��}�C5�)sSVe0^x��xN��d�Y��G�����=ME+BY�$��`%9ǎ����ol@�-VΡ�5rJ�����J�ڞ��O�zqm(B��C�xǜ̃%�P���O>e#K�KV6�>	mG�I��u�L�&�R�6 Ҟ,���Zhd�\�-k'��˛{�K�X���(�DhZ&y�ĳt�^G�o��.
�^uh��y\IIKRTذ�)!;�^�"?�J�ߖ�zs���F�\�$��J�4�ܰ�ݏ��l��,sY��S\�cfԳW;]�'���!���4,b�a��`�6�MSNw���p�q��#�a�kJ�p[���YLw~Gī���O��F5�Vn�0(��(ƬsW�Whd�S�w��|�'Dǖ�K,�Se�ߜu�"ɛ�o�(�q�HIO��d9H*�D;%��,�UV�")����Ν1c?7�/��TֽJ��K0���0=�t7��w�}I��,	dT�)�X{���݉��ͭ��Bu�'"��X�Rܶ�b�m��k�N��O�ʘ�|\`�9��'�hg����V7��(F�cԆ�χ�>0Z��v��[�c+=�c	%�p�����@�O�E��nH��!�G�h�X6��k�rXH�	�3L����N℀�k��ϖ�ۮa��Y ������EZ��G
$����/Ez�|=��K�2����}�"i�M0�X���-�$�V0��g�qIg�p��pEX�#m�:9���WU\V�V����読��i�?dI�[�R�����c�h�"����(�_ķ�\Y�gW���
�qq�m�6�����v^�D�ۊ�%q��.(�7����M_y��P��ZC����������{�n��7���:6�!v"�r�gr�Ԙ b��L݋�n�K����\�E���c���ε���+����ރ��ȄN+����[�����y�yK�=����d�oNE��h�^�M�8S^��8���ia�_��j��1��G�ܛݜez�0}qW���S�6�{����̯��c��n���������g�9�?~^��E�$Dҿ�N�HQ8�������@��z��3�B?x�p���2�-��T"��np�O3V�9��M���!��;N�T��\"A�Jl����������)�u��v��^6���_b�y�o
/+i��u�L; ,�g��h��傶�+�YR�I�k��<#{�}Q�3�aiy��Ϋ]���U������Y5��<�}�Qw����2�[)��DD0�$�б���'�p1�]�X*��>�8)w-,�+��Ya݇S�Jc�1��d��§"���]�ԗ�+o���ߪǾ�}�{��Е��E�� �xـ���k�V����k�9+�T���RƊ�S��\����f.�DIW����(M.���S��C����>F�p�Ł��������.u���b��@f �={����#6¡���&�('�|�͕��BI�k���R
P��羄����Sr��W�n�X�<XA��)���������������z�e� �\��&d�p��\��w�����p��_�Q��OI���tO�c����I2D������D�O"���c'y��c�C��_���)���G��� F[q͂���xKn���@6�fiO��f�Q����L7r#s�jf[�g;����tk���{�k�<���$D�;��&�s�TǷ_�u�0bЋZ��PnXY�*�~��n���3�T.${V&�R26r�B���ʖm)03���9�\<'N���i��{����u�yJ��Tp�Y��.�Eܐ�Z���!s�VV��/)S�e������Gw_��Z��J��X�8%q����(נ-�+��{�%]k�-�%�ү���������m�Mk�9Â(�;���õ�s����8��E)��P�t)փ�<�dE[�}G,/���<U���F��̴���=�[�:��UY}��m�Dp,��ioPC`t_�)z�T��=P�d���Y�4�\5�%ofh� 8 ���.��}Kl����<g�C��d�C�<= �lc;a�G��	���#P�~��x�C؏�_�ywq�d;$���tw��DPPK��#�X�6[Rp����d�.�Œ�X?ET�#����a�l$]]�Et�[��te!{)8?,�(L��p�tm�{7�Do�gk[R�.���ŗ�T�%l�
��8��֎cӗ^�FZc�)F�үd)k�̓�n��HP���,s���o֠�\����D��TK۴�Y��2�x�tt�m_'���EI� ��&��F��%�hx'.������eT"`����&2�����Lu���[0�˹���;7�������B+�D�{���IT�|�������.�	9$��F1��הC�-IWR�(��$m+�j�ӭ*��ď�&��y\[Ġ3a�3=Gљ�N ��S���>֚s)�k���O���2�QP�|=�z<HRPP/Jʜw/+��e��ߐ�Nv�6�Ai[(�2W^���5�:+M��>g�JtS(�o�<�P���`�|����s���C@��[��f^Iq{��ھ)B��C{�c) �qE���>�s�W�@Z���=�\���u��$O+���9SS;��f9&<�
դ��\�\+��=(���:y�^.W�������k�!ڡ���l`�$�5�k�m2�z=q�C��e�$�b;X�`���lj�}��zG	_B�m:uҩ�~�$����]+xY~��r'�{��D�[\���؀F��&"�K���so��)�N2�K��L�%/3�LD��b�B��_�[��;#Ʌ
���zg�G���m/��<�{��kY��mQ'���^�|�
�k�?�:P�T�����/w7���N�t��n;�LB�LK�VX���u�#-�ZQ-��'r�_�Ȳ *>��;����S*X�3:�+X�o��C+��C��W��=���s��T��$��{�FV�Rd�N��;�hy��m��ܖ"�f2��\�k���k
�h�ۍ*�M�IG���Qƛ��X���w���M�����dg�l%2?�L����ŧ�Uh��ab<��r��24����_�!�u�Z���po"Z�� 4��m^��qd�qS��b�C�i��f�2���-�ƒA�}��q�d��.X�E�a�����_�ܱL�6�uL�!��@�!O�a�j�"��� �5����ڦ�������"<eA](�
�JE7ǉoߒ�~�w�p\��+O���W��J���\��j����u�U��,7�Fk�ɼf�YoCkK^���X۪6����*�������u�^��3�Q�`l�~|�,|����M��v��0r]��TzY����^����KY��C������/ug_���_x��h�9��:U��LתĶ��C%�w��1
�ɚ
�F�}D���qC��;h�+hG�����J��Ιךkj�������b��'R�&�/��Jω<0�3֦S;^sZ�O��LU�xt�]���V�uO#%��ǫ-���LjlK��)=��[Mu�����N%��Jz&��ؽ淫"7\�-x���z!P�~��󉽑�-9����S]�_�f٪K�vAu��Ϳ)i����l멗!�2,�P��3��"��i�c��r�ˎc��q���EM���y	"�~  �a4ngᴶJ��66�(D�3�O�e��NY��k%�٤Ԓ%�����^��+�*
B����1��qu�����e!/�~��x��1���q�Vt��47l�q<�r�k�XT.%��1�%>&�U˞��z�����Uy��k4W��Pv&b?��&kY�[e����,Z6S�},��W���\��<
=\����r��U+}�v��;�
�x(��p�ȑ=�M̑'p�чr�w %�s�:_(�N��܈�n�H_a���Q�2B���q&,�S^�R
�%u_Ņ���_��H�>b_)]��J�NU��*yZ���eDN%�HwO/�N���a8(f���WIc���ڽo�Y�y��:��}�?�g}��#P�����3�@� ���3�-���Ζ�".(���SB�K�M�5$~O�a��F�[�9���cWx�c��c�I��7
�D��ͅ�g*9'N�Wj�c�!5���뜒���^���Q8ώ�I����g$m�lJ�%��/��hw�<+Ơ�VوC.�-I]��*�l��w	r�=o/E�u�/9��vץ@����ϯ�ydK���������t���p�S"�%[�O�iZ}��|�O��M���V�i�3j�������s禮a���PF�>9S;n�uN���w\���mpr���R^�"I-����v%��*�iT���r�Ż�tY�TěB҃��Ϳ��Ϥ;O��B�N��R1��KEΞ$�d��yn����h<��]c�ݔ�!I֑�O+�wbYS>/�Z���^�oU�ޥ��u]]?�X�p�^�A�;�ݞMݏ��TMA�ӗ��􂵱�X�WƫH�����?����G�����bc��ˠ���}��ά&`dN���mMN��p��K�(����E�'<Iނ�,D���A�,�ɕ��p�Ҕ$��>�w-ho�D��<���v	C�i��n\("�ZϢ;'v�JBC�Hb޹�Cx�7"^��V��-��A�*L�=W�\��c�Mu�Ľ�,?[��e�ͅ-&�sM���p�A�8�^��z�r�n����[�]���}i��yV
�۝�d_)��?���PԤ�tS�ˍ���	��h{���RP���֥�Y�{���+%(�oh�w�Y��+�Q2`i�o"�a�d�����̧��R����>6��zi�p)����f�#
^�(Ir-O��ay7{���m�[��<��e'1��e����I��zl�`jn4^�lf��]�^�e�'k��	)Y3�ϹV-LTH�y[�/ʥ��4"ᐬ�T�vI�A�{���*9����%�yކ7�㏲��@[�*Bk�"I�.>co�ީ��0׋$�^����@#.���8�P��A��p�;�9�R�w��5�����5������bW}cvܐ��n0f���Ԁ�(&{�������ܿ�?URS��#�'q[Z�g�ܗp�F��<�WZ�{! �Î�[��߃��M?LR�,/��mV�ƕ���{Z�5��V1Y'���
QxQZZ� i��Pt�(H�?���;��"���k-�L�5c�u�Q	�����I毽*a�ԅ�h��h�x��J$<&;��RV�1o�r��31ѹ������n��qxe�߽�-� �x�mm��d8Y��A����)d�C��3��N��� ���3Ͽ�P�l?�?&j(Gm%F��d�K8�8W����ǲn54�(�3��²>� �ؿ2���2�슧�$(��hW�f�gX���X��1�!�Hy�}���������O{�l��짛���T�V�sy!/�IfN�� P���ԧ�L�C_�w��G� ��	�[[�D�dצk��a5�l�`_������I���i���1ɢ�ֻ��]C�)v�Qŉ��G�Vt��]Wx�Vw�l�6D��a9]��aF<7V���R2>�@Y�]�[Z��>4� 
�Ɫ��Ȥ_K����S�q�S�,�����&3\�˼��d�� c���q��m���JU�Q�.j�����c��˾�S�Q�X�8:��#����$\�ky�|f}_�u�[O����ts��\���>@��6�L�ܹy������w��:����A��M� >��Z� ��P`\8)���2�I�7�k#u�4��AEu�xf��X>��l�c���DcB�Yj�r���!�}n���0d?2��<�zV�T^C1��ꈜ��!v��T-����V��_��|rg�ْ�X��������re��X�E��ݑk�Q�z$1��r#t�t
����xv��+]��<�^")����K�t_�˄sv�\�)Ȣ�Fx����q�'�h��QD�X�S�5���5��<'mYNYP}O%5����Y��HlВ�@[���5���diG��P����?���\F�'�ƀ�%m >^S�oK������^[K�F(0l��5�]�L˹6�-�'�|L�^��e;E�C9�/d���F�`.A����uo�c�d����#��)ƹ�F(E�W��~9�^iI�g+Z�C�/�Hi�|]�W^�V^U��:my;��2�r5���J8����j���Ś��Ã�~h�q߾�A�O�wǆ�>����!�NG.^>7��f�I|��R�>��?���Ͷ6�k�]��ɓDJ|g�� �m��-P��z��׋�Y!Nz���>���B\�BH�W3�Y�Y�~Ƞ�~��^����K�����a�����w�|hݵ���v��>��Mșxg��CBX�X{�XB�g�%�,t�C�����K�l�����Cp¿�}���u���W��<�Òu��m���N�
,���5����w2���q��vI���<-'S�����^V0X����L!r��r1�v�1I��oCQ�$��Jv�Y_d�E��a�;�3{zД�!�{�ZtϞc��}�x�wC��:!/�tC�$Y���;6�QaEA�F)�C	~$/�����[�]D&P�zKR��n��˳?�o�<B7�ǠO�_�$�_s�~oDv���#�Пۡ������du�]B�o���]q xB:���T&3aA���.��5K��j�B�����.��UCBy��<ߍl�����݌�0���"���v�]�q@��@���Ck�q˨̆�;b�A~�?�%���DX)Q3E$2�y�����H�)D(
��&1��u���k�C��mF��։Ra	f���⏬�{N�b��=���S=㳔����y#�¤V��b޶w�C���i���l(s$u�l��� aښ���Ӯ�ɱ��vS��� �����4�K?Ԙ�%T��O}B�(I��w�4m�iT�֧�]��P\�d��)q.�o�8��#Z�H�ñ����J��j�;TZ�=	����a�?�޲�ЍǏ�,B�͚k������K� 6gɯ�xn�tE[X��L!�D����e2��>F��΂
�����ʰ�C Ǟ�!8mq9F�'V�t�w��9c�hCq������扼A��z��o�0K�dGHq/�Wm�Z����9�A1�ȑ�:��4����k��M���8�$���X���^-`����9��PqJ
L�pf�vps���Y��ŇqlZ��=Hb��(�Joq��K��@9a�3��yg/��Y	���A`ӓ�������!I�s����G ���y*�M�H7{����4I�,O넆6��Q�O�Q�n�V�X��p��3ù���ޫ���0�#C���-V���H2g,�w�����8"�X6p����-�"5��]ڜSs�0P��s�|��k��M��uD��:��}���oھ�Me�#	}pn�*����oFM��约x�o��s�CkŮf��E�Uu=,�I8�i6���!o`�m�l��IW|o��v�:&�䳾�G��d6�/����3�"��di��E�b�x��B���d9Y/MR?������+X�f���&��-|��[�C���uS�~:��8"z50�v����6��#��aJ�!��8���qq�P�R�9Qa��p&���W��}g��c�����>��L�mmL7�����P11�>,��	D�M3w|�0BS����Y,%���ys�7��{�A?�\�����M������z�B����F}Ҳ����՛k�@�5�'uGB�Q5��!h��'CXĮN!�v�� �^��{u?y�5�6�?�F�'xZ0!z��g��6�>�_�Ԕ��-��!���I����X�?�N�(�l���Ԅl���7x}Wd��r�]�i��
�k"SI�����}�\ϫ	�J���4b
�{(MA�W�v�e�2:��� ��Jy��a�:I�3���H���<�C���e(V>\@(w�k�y�C=i��z��7����}X���}����W�=��C���I��R�1�����iw��KK�-&�9��]d)�m�n�a�w8���u��+��}>C��nxM�t�V������f˳ܰ�y(BF�Sl#1�ᒮ��HA�����u W�X:e��$�pק9j��H��g�Z�8n�V`�L�J��,�
b�u�M0B8�%��$�$�^Qi������$�yng�����}O�a�3�Jc0ER�"V6���I�un��Վ�w
C{�+8I1K�f�#9-��m��ч���ǲ��T$#��q@q���P�rM���p�7/��#��\qP_���{ 1�X�9wbpsN�e��qky|���X�o7�+��Ŀ��n΀$۶�Mx*�2H�6͕��� t�&N�Ê�#���{����3L2u�@�T�T���>9'sޅ�N�I:���ʱ�;s���|�F:cߊ��D�L�c2+�� P��r��T��S����=�K#��ϲ�$ED�&R��ֹ�~rTs��>�2��or��)����k^q-[W�����L>B���9�:ol~hD;�;Rm�X{$��v-�]?�dת���LV��������;å���^�+�qs��C!y{䱉���� �FLQB�����K>�<�7N��Z��9� ��<�"�x���ZmUQ	xc�W#�Ǽ�甇,H�ag���Ť��Z�q�rc�X,��O��b8��Y��[F���_���pN������v�ሡ��}E\�y�"��gY���~��c�{�خ�;�g����)���#�񥹯ڵ�����0�	�/���T�>��?����6yr�<m�7��u,_C��+�jXr./i��<+��R�<��,"V.B9}�{/�w�I�AK�ݱ�T�7����h�?N�H�N��6=�A;L�Y+��H�ʋ�u>Dݷo ����߻��K��ҭ���Wp��6�,���*u�ܝ�5�b��	o�t5������"��7���l|���S��ϳM�A��x�{/�����{�N[{Q��_������*�h��QS:Zs��z��_B	�,�H�sb�{��~�)��9�+�1�ʓ�p='r�@�������9�@(0��r�%��9��	�t���f�s�6�vq%���G9?���8�\(���.W�Ja(�����!�C#����G���D��v��z��~1�C��@������zu�-�T�}���]���m������%���\	kMH�W^���)�:L*�;BJ�	�+�ˤ���R��@�Tm�C(Q���1q�W	�k,[d�L�-;�#D�vs�Hvh��Gk�Hi瑜��Lnj��5h�����Y~��$�N�����a|�gX�ոg����c����%��C��~�U�+�`-+�-�)��f7wTr������vM�qm������%nm�p���O�6��u.�㴞���:N�GÄ��Û��4%ʟ5؛g��eȃ���!&���ѽ���N��ij\�s�5���
A{N���w#��m�f8�����a�����M��\O�jBzٵ�_�!�u�b� "ԋHZ��V �>[Yb��;�DZ~[7li�q:�lI_�2N)����tQ���1��3�
aCRw��Oii	��B)�k�D@�!���v��Ħ�����;�#���o�[zm��q��$���6ln�5wp����Vp�5۬�TT���-�ܨ��@���x%���A���9��5v�f�Z�@29�n�Iv �J��������1i4i0�vd	D��:�C�	�/��;.|�s���KbԦOL���ɩ��V@s�4��jM9��Q\[�_���`1N� �h��w;���DMi���?x<vV����\�:o,E�����mM/�����!��Ĵ>���m��v�>��_�A|�.lG�K=W�?�(F
r��7����edKbr���0�}NX'v�Z�2|C��jq��N5�'*��;��Ma��wm�p^�֋�9%	�R��F~�:b������a���gQv5�SS87�qS{���u����Dyp�SI�p��vF��E;�>����x���2����n���euy�����&A�����|� �t�{����Lh�C�	-�%�ɘ_�3ٷ+��D��q���}>R����6��	iN6:/�?}[�^��W2�R���n�>���^��/���q�9je`�O����.�c�s߉�a�DK"cH"�Q�V���n�_�}B���]&f�Ƌ�a}�$�&��:\PU���'��#�l���`g�H1���b�o��N�Pb��;+T��b�Qy-$�-Lb�Yj�#4݇p����޺���&�۲�!Tk�G�����z���n�]�����3�Iy���V]c���T�������Z�y�f���e�ϊP޺Ş�l�4ͳ���ǕP⬅ᡉ�;�����`r�-�����5��b��"��~�zv_��N��@)F
����i^�F�Cr���9���j���iińC��~F�ۜ�O�c����tD�.�����w��<7��u���'��r�78HNu�`zlGo���P$<v�)�N�F7^ua�K��P�g�e��6e���\�G���]��م�;*�l���O�Q\�����a�(3AK��x���B�Z�+�;9Md� ��z�`Bhy��e6�J��d�3�K
k��|��-�9eE;+��xӓ�)޻SM���jjI��.��fb�ue���K�)����$6�/����(�Vc�2�N٫�Ӷ}���o�/lO�ajˉ���Qz�Mcq���?}n�n\"��V6�~�����ջ�^���Y�
��ݽ�;�)i���A��`�]6�u����
V"B9��1 �&j�1���ʱ� AnO;\�(U�!\ϵ�������
W�82G�"77�X	@�
�-�/�*:���V�3�3me�2�VB�r�3��.���:�%i�]v�q�����\w&;������1�t��'f�&a=^��_�a�N.�#��zg>�mb�4��A���X�d����VZľwV_� =ҕhb�&LTo%i���jB&����^��NJ��M�-PAn;1�l*�%+������X-M8� �e;E!ܠ�.��n#�����B��A|鈎6Xp&e?zKPrMs�d�A����=���c{M����a2I�����$�F�|L{Vd=�$�El�fbS c)Z(��<����~�X�k/@��Z{��O���+|��T�bZ���������`_�"r	���j��3:}���o�¬���ڳ��9��9H�E/��a�f3d�[����k�2mQ���$�Q��D�Wlv�9��,?9G��ᛲa2W��[�߯W4��0�ε۟7���V����U���" P��"�r�q=�,��ٯL�'�F7o�S�r;_d���{Y�,}�+�2J���m-[�����'���zMA��4t��aAPC˻e���}��P���*#z���BjM6��5)�%I���B>	KWC�iDE�hbX�d SYk��0�s\�k�P����e�2�.�|6��[$�͕L�w{���Ir�P_�v#��\N#Ɖ�����)���i�G���+H�(�T��4W�"xY;��s%H�s���#�2��a��p����Y�v�K=f#��̷�bl��msrgb�A�4�9�W����~l�J�C���g(0���#��~IB���$�Fz��ބh�>�U���}�X���_lYc� ��۝��L����c��w[�S���@!�(�L!CW.��o��.B�ƃ{ص�Ǐ]��S�������8��4zm�iW1�^D�m#���HEϵwsU\y��3����m���N�8d��[
[܆���}�B8�1��֊ݳ��(��J˘����Y
tNV�R�
H/�C~7+9�$M2ܛ&��5mg�P�>��]��VO�bw��Odڔ���Vr��E��2�uB��7�'�lbˈo
�p�cߔ� .�E�������$!�P=LBI�a1�5b2�B�����΄��s!�a0`���m��%�a,�~�4\<��#�	BO���4�Ąb^��7O�U�<Ν�7��E�#���J���~bd{���A��o*q�����PJ�u$���>*�*�:7R�oJVv"�.U�Aɖ������g'���۰=���H�p���b����"��=������W���.W�76s	Gy�D�O��F��	�asY�T�RE0'�$96�̈́�[�I�M�FP���l����D�G#�a����
�ic�$��2�u{�ڱ������CZ]wI"_���2Ԃ���5���t�'��O�B�D�룱�����%�^��-�����q0x	=8g'�m�'�5e�g6Bm�i��`ԍI���3�%s^S 
�0ё�m��Y<�_�Ɠ��G:I�"��{[���e�?��mLq9'^}�<��'y/+c�c�=t���91�K����2*M���5e����R��m򽬸���w�ư)"͋�\�1*�pH��n�#gPf_q��}f/����G��k��l��G��[^��#E��qT�Ч�t��j:y_�?�]"N4S��XW�KO����2�߅�����߈��ӂ�s���������kpCGY��g�2�{"K7��f��v!�e�8^	a��-y���,�$@�����5$����tG��I�c���M�6g�q#ڼ��Ek���>��z4���$�F4�:��$��<����o�\���jB'Qpge;РP(�>�8��2�&�$>��h-�)��I�]>�^)hnv+r��IW�-�AB^�iG�#B��{ a��շ/`t56�����{�	%�]=�&YQ��wއ֯�Y�^+\&f��t+=y]^{eX(��[
�0W�r�r��� ��;>�Z�]ڔ��noZ�(�X�<J������`�z�!�q=	y t�b���㺿*B��#|п�����h��h�d(
�X~B�d����;ͽjK>��z��$u��I�!��ϫ�~hQf���В��|�t��^z�֩��8�憰l�$��k�i�/�Ѕ� H{wm+ ø���\tb�;�m���7�Sv�J��͍_��OA���W4V���^S	�Y��BKM�|�;���	>L�Td���G�j�2歠K�X�i�c�+	-�:��Z�!�$��;����]�YW-,�9�;"K5H:��q4>џ�X�d$e�"��#L���3ٱ��s�c�7G�@('�Z�{no%'���v?�Ⱦ�v��ZhEe�q�+/��E��V�֩$@F��==�XI�b�Y+�y�#q&!�aԬ�V��eݣ�{�vb���S?�:/�����#P�~��X����֣�oO��X~^���]d������g�C��h1�D�Ln��/C���oD$��*�tD
�hLB�&�ޅ�!ՄoKRj��v��i���iC�a:�y�u��t�[�l@�.�j��-�y�fσzBiD�Mp~9m� O�6Sy�Y���޾C����Л+>؅��P�R0Yӷ �!�n�B�Lo�3O!��9^&�������|m�����9a���Ƒc��)�@�ydx���1�ܙ\��^~?�������������Ƌ2�u�f�{{5�@����~�<��c�\�7�Fn��vd�6�c�[�m����{��n��M����D�h.�D��ѡ���	Ӆ\�Tl�O��qw��̊�����o�Я�����Ɠ��śr8H7�AK?��	"rS���\-��6M�Vb�ݖe+���F�rī�g�P�k�df���2����ު��L�El�e�,��0�V�]�nJ|֔�a�׫�J�G���0��htݾ���M�I<n�zI�[��AX��Z;E�8�F�sp��<�~HJ�e�ڼ0}k���\	�>�m�h����^�5�b��b�w7A#���������6��5���r3�9v�0g�֯]�D`:�k���)7�N�*b�����o��ƻ\����x��C���N�܉��y1�l��l��7t]��_ב��_�х���Z���ِ|�`������Bp�6���]e(�v�>A=�Ch�lEt2�>qXE�YE����6����-\�:�]�I��$�oP "\{D�G���v������;��c��J�ՙ.���E�p��v.�i�Ν^9<�\[����O�']��йްhNO�o��G�$8���6%,������mK�����T�}
E��ʮ���@��v����ëc�k�П��������g�!5���ҳد;c�X�f�w@��2�g.����֚&�F�|�D"XBq/�� ~~(x-�l�d�R[���g��D֫-�'!=��1�;f����c8���9u�<���)?���1��w�;����]뭩C�*���ew�t�%=1{c��ʇc8��V�q�3������y7�v�&�����[�S���Cedx�F�v�F�yj��/͜=K/ּe(M:��o��р����R�턚���58Z_��"�e����L>�,��_��8Z���~�=�X�����	�
��Jk�`\B�ꙙؽ�%��5��<�>��]��t;a�l�<���\�$	}�D�t���Mҩ6�w��6`ߝ�w%��1�lw�X��D>$�!�G��n�ݱ�ڹCo�!A��8p]_�������^�q̢ߛ�G�.G�pnF *0�}��c��O����NyK��p��{��M�A�v������{fI7{�r�g4�i?�O:5���(E�с��6k2�X��C�B��z�<b��b�&c}�j~(|�_e�-����{��Y1�c]��0,�4o{맑� *��n̸�17���c(���O㗧)/q�.}�\-�q�L({��PK׫-�a~B���k�3����ǈ-�?�ז5��9��n���ޡ�;{��w_��L^E]C7yã]�i�2���~�^�ڷ�ј���p?��\;����f{l����:����X�v���o��y*2���E�O�_��Я�`>kWT.w��(��B��\���+���⶛/�R��A�]�;�9��G���Mݗv�����O�� ɰ=C����h>��*�c؎V�e��Udwl����w�J[�p�r�z˰vS�na�і�����ȠV�=�,�?Tbv.�F�;+vwl�
��p����(��WqKk��w��\�`7N9��y+����=���y��O�65Ʃ��ȴ����έ�s�%|@�g$�i�(�~%�'k�)�/; z��{$����@�����^�Go����n�nj
��C�zH>���qa�˧���0*~Wk�Xmh6�(�ϥJ��tg=�´�+��4�e�T���!)��j��]�{�mg����kb�Q:�� �k�=������C<ZsU��Y��ƫ}��o�MVm�X����v����mhY`;%c<���?���w�v}�H#;.9���E�<6
��k�s���Q<'/H���(�t��.gYb�����gid�\!P��\ק���tr��9�R|N��u�)[�$���6K�f6��gyR��� ��<��!ɣ)Wa�xhU���d��vSZ�����U��P!jG���Л5�^�t�'a��mO���_��q 1" �RSB@Ri���M��Ĥ$� ���aԂ��{����?𻞼�_�u�����sN�;F����� ��0�O<7d���� ~�����û�||k-_�C���<f�U-�B��q�W6 ���YP��#��*����§�/����m��> >�\
�"{ci����]��Y����5t���0+.1퉣N��ڭ�X�N�\�Q���k\��Xn�__��k�:�|�?����C�g�&�Y�d�/@� 1�C��t���>��������e�oD��?VD����g���$n��j��s��M?����N(�f��#㚶~�� [��NN[�0ς���z�sU���*\�f��|R�ˆx�ٌR��mɂkF��7�s�{�Į�������J}^����_��UO�@&�|������Yx���޿�j"��)��`4=4�������<U�y���a��ܸ[`��f����R�kfe�7��\�8� #��S=��OO3�3�?S���M94dT�:���/љa���k}E����FjW��%������_Ζ�9rCv�6Q3��Q�%�b�6����K��ݕ�
��US�?w�{��~��kKf"P�V��5��_���g�	?���Z�.S�G*6,����,-�D������4���y,�^����u8BJ��_M�2	�Ձ{T�ʜ�s|ݤ����*�3�S��B��.B6��V�*4x��6�W���Uگ���5ÖL���R||�J�:���oſ�O��%G+���XWY����v{��o#�6Җ�rz���l�.��E��D�$��������<h}�gb?y�BΘ�1;y�0C���ĥ�e\�.1$�h�W�_P.)�[�Ǉi�OG����o<�X��u�X�A�Y����΍\�6]�������/P�g�r�	�jT��{Gi'uw�]R���2���B~1������2��|h�ݛ�俉|K������*b#������ox�U�c#@����Ҕ[�n����[�Gs�K\M�O^V�U�x2c���S��ET�.�����͙��+֚ŝm�W�7�@��3���;գ=+e6� ��F#�uE�i�xM��k�{�?Gb�1�(���흎�[���>~h�w���{���)} #R`2Jlt���`]C�K�M\v��g:�}���������3�T�"�B��=Z��v�����ߴx 9Zx�ͨ�JZN���A�8M�]��Fx
���Gab���yf������!��d4
~��Aw�Z��O�\��yUj{���ީf�̿U{h�t�����(�!|=-�;�&?�d�����/�kZ�X�[÷ IQ>�$6�񝮢:�ܔ���.���R��p�Y�����ҋ�@^�-{<v��er!$H=����z�[?C��p��^���c�z�^��YH6�L��}�+G���Lr#e4ކLl$C�S���ɖ��3D�=N�x�����E:�ẝX�h��Y�����E�RV�|��^��<e�u���Qj�IKƱU���`@���U�IE>@yG��Jk� ��٥}U&-�{x�JT��߶�����^"sc��Oθ+t��xo������{�l[�A��G���dl���#)`��»_�.�Lw�!S�t&-5�匏|�w��.cش.���ᙘy\�n�x3z��H1���A�i��z�����]���D�{AxX�L�]w�F:]�n��<XW���Xm��c¬d�ظ�D9��TƷ4���'�������aM0i�!��.�1��"�1Sq��v�;#�!m����]�#]�z�Poϥ�Yw��P��#�ɭHk�=Č/M�C�u~���q�ք�z� �4��r{UR���t���}�(~�+*�c[��n��|(d���Hn�=�s��z7��͗���c�z�Uz�/���kƄƥ9r���s��`�@�˪'���.�+;u~W���̯<.���w<���S$��)����3	�;�Q���t�Rb�_?"��${d�E�tG�ς\��Ck�|X���Q֬�j���s��y�����-ba�����r7�����&J�F91���j�ܟ~�� ^���%�ձ<Cf�ֹ֩&��i�D��iXs���Z	��$�s��kf���R­�*�f��0�|�޻�ek����BhI���:�n�GA[�\�,I��ն��~~������ۭ˛�0�����ހ\Ж���I��\Ǎ<v]�~H�>M�d��.!;kK/qxa�/ћ�(j}P�а�HG�^����L�ʟ���̂%^��l�.�Gx���������氰�#L��ȩ��"ԛ��:�p��' ��	1k�m�v���}f���-QJ�+�u�+�Nm���_���ߏ!�&�p���~)wUb&�q���	k�u��N�G���x��^�7�C�O?�a�
K� ��3���:��o�A�����j[\���>�/�xx���C2y�m ��%�<��%GwA���愮$��#�u��T������{n�36� � �\%�k.J�y��f͵��o�l7�P��,D���Uu��	P�w�t�\���t�s�ᢿ	����pD�}8������m'�-�$zCu��ُ�سr��"��ؾ�঴�������}g�����is>��#CI��ÒKBrٔ��=ً�r����]b�ѣ>a�i�� �KNʺ���>W�02G��2N�8��;���G���?���t$J_�f�3V�4�I+)	\�)@�wzq/���<�5�h����V��5�l=�*8I%�_%Ȯ�pˑb ���~���K��J'��+��8�����/RP?:�RzZ����G��ڼ;�S;iUw�� �+�;�`�c�2�Bǽʠ�� �e��K�t�t��Ygk��ɯ?K���px�����^az�7ｧ�3��~�^�  Ks�z�uM" �5��]͖ؽ����t�֍ KE���u���/���m�b�'͑�=0�����W-W"�A΀�i��F�+=ы�4�Gm��5��GĲ&}���lgN�֢�6;�;��{wTN�)!�@����*�K��J ���),�Du��.�S�I���6���0��a���NG�'��Tm惯��O,Ϯ�DPGb���K<��`j��Y�
u>�'ڕ<�Н{o�Zwܔw���1��v3;�^:nv�*5�bX�چ{)����@ߏF^3
;goz���Bn�|����^@�QW%ӕK���p�B-kWۑ%�(g�������L-�\ɩ�"�q�P��
&��kPM�ag�ͻ��)>���Τew�/SՄD�љ�qvgO������ɬ��szeϾ��/��p��BLZ�/���4�}V�z�p���"�/�����|�d�'���|o�#���7E�x{V����s�
�&�d�g��&���G�����O�W:�zkn+3f�a	Y7�mݖ�zZ�t�����/�x�Z��wK*>^Ow]&=_"��= /.lk���~�#�?���T�=����ӡ?�MbH���t�I��o⏥�*Б,7�Y;������D���cc$�Ͷb�%H~|w?���:���D����Y'>Sݵ��Az���e��ȩS������:3��g�e�ah3��P�yu51&�Y��[���]�o�`�j�mD�]�/��$Ot�S,
������0��`O�lQr���)��KSՊO���<5�^�������r��Rl�GzƘ�]�k��&#��٩*LI�h����x��Aע��xG�d]@�%�E����̻�v��>w��T�C#�̿PL���&�eϔ%#��c6N���C��@s�d����S��Z����3��{	2���gne7~�x���g���>5�˟���VW��}�pCI�'��LtV��Z��A׾w���r$�.����z�,c-�h��B���i(6ϣثbW�O0�`�h��[e���U�EE�tp�æ/�}���]3�TT�VmZ\S찖�	�����ޢ�����g��A�����8'm��S�#�Ė&�:�\;cx&�������α������~¸�S��FqL%+?m���Wv}n���nф��Ev�3(?����mٵ/U04*��]�}��U�z@rLHus\�Z�	�U���tױ�a�q���7�O|�^&W�3�En|��Q�.ү��P:w��Ʉk��>Uf�z�,���v֤�AӲBN�%�`�9��y.�+�\�~���Л��%�!~���ƴ������~,�Y��R�*?@�(8����-���?UA��U����٫�d���L��U+}�^�ރ]Q��%^�Y��W1X��������0{����K�,*��<�ׁ�(þ���i�{�Vԡ����2=���!�Ɇ���>Ƽ?�(�����@�˄:}�&%1jI�w��Us�;Тμ�zl����o\�H����Yw�#%ʫ����(�;�oċ.bʕX�C#M�����zM�/�Buo��,/,�������/��������9�������7�uWUI��E���+U?��mؐ�Q'"X+��K�`#.%j8a��Mi�:/����Q?ʈ6<7�3W'�)�>o�"��޸�qlt�q�k��X5/���X���Vs�ɽ��p�'V��Bѿ$����)�Ġ���QsU�l����~���@�V[�|j�s�����b�t
����>�����B-nE�P���a1�Ie����c�����!y@/��[�[
ɲ����	ݎ��a�߉n|n�z�8�~����*ت)-w$[���e���@B���t�5o>=~ɓ �f>�1��P�/��T *-�����r�m].��t���=з
U�M�
s����>i�ƺ���אx6�F.����2�y_�txM��Z��C�E�hI�V�v�*R�ƶ������������ay��ox���T2E;��Eq'7#����}H�f$��I����U�am�����8�]F)k��[t�%�=�n!�[4��-^�=�ϼ�z;:ӕ5fQ>lxY&� �} j*A�~��Pj�u˘Nq��j�H���i�'��u�z�������nf(�h���E��h��)���8���<bb*����L���|g�1Ycr[|�{綻7����?�e�>�������Q���(vO8�S�G�d���s���X�MeW��,o�W)n?�	�S=��a�=c��BtWd(t*�t�u��ynd^�\.;�s҂�&�V����Eo2��C��3�g�+ �e�r�1�}����t��i��䌟x1�5)�8U��T䃼/�� l���M�n�NOD9�mRw��q¶�^؏����#��WM8KMQu�G.��{��N�>]��3M�<�r*�<��)�0���{�'C+���T��ܽX�o�%Z
�_s��������¬�d�_��ېÌ�o�ɦ��r�z �
�̐��g��Ղ�N�b>Y�o�8��K,0e� `�*t�鉠�
}�S*��%��'�vJ8Y�����/�b�'&��A���7ܹ-]���m���#Ѫ�3�s��W�fo;#v=ϭ�2փ5�nr�}�IU�M�)ҭQ�iC��`�csH��h�?6�I�a��QPV������C�J���]�g�L)M�����ڪŶ�����v2��)� M3�I/����CMۉ�ŏF6�&��T�m`V���Qx
}
����M��)�i�<�i���W��cd���tOV��sS�Q�L�	�S''�<��f�w&l�kZ�`V�ً�r��W=i�u�^���Q��Ƒm�������G���-!mmc��c煓�E^����7wZ�5��X��V4�{Fy�~��I,������"ʍ��6�+�&�v�X鯿4��2)��s%��X�5��4�2)�s��V��e˧-�TܙY1�a��$�4Cj����w��w|l��&!L,��0�M�����C5�:,O���?���f����V��~#�ǣ�M�� f�S���Yc@����2�*h��̆Fp���V
 ڥ���)#Jޭ����h�uPD�&U�;\b|?�C~�U@�����EG"�S�g�Ě�^����Ow��C:�f~�&L�Ob���	{[���ЭB�%y����Y�����f������Ӡ;H��A9��j>Ҝ;���nⲩ����9�I�{�1��/��� ��լ���9zV�YƁ�U��h�7lW�Z��î������9g�ǅS� .��$�R% 4G�\�c��_�n L�,�6��%5R��ʶ��C�����-H�Fa��Tf�Ҕ�<��yjO/�§���N�3��GA�v��o�h��ؼ�WB����ld]Ó�a� X�=���Z25%��v#Md����Ql�}*>��\d�\�_t��8c�����#1Ձ�vq��3��d,2������Jv�������Dli]�$��?�z�`w�Ḱ����o	ݑE�S>>A`���4�LW�A>ֶ_���v8U��zo�'e�aJ6�f��AM�D;�~������N4sR� Uz��ta_�(Y8��i$������]F��*��
C��S�bJ橹5�3B���O�Tս�R�~�}��gi�+Ÿ�=\��\�H�ndL��5�x��.BA��u��� ..��}!��5���S8��b×��Q�4�^��4�}OH^軣�����������w�0�y7��Ԍ�����˓&Y�83�8i�0�#��y�s\����1
���ϕ+0ig6GG$~�S���6;N��2�C��^�&Aq@*ma*6z�o@Q�0X�n�$;bOc��A�b���G������O� 
E8� Oa��8-NZ���@�4	H�z���6Fz��]��?�mlt��H_n*g�H���4\��68�/Sf�w_в�U'ȅ��U+	��Y��?6/��S���� �R|b_���mj����UKoN3϶� � �zF"�=]:! ���*�<��J��ic�D�'��'���'/�춖&�íB�jMʠVR�91��Q�]��k�!v�9�mY��G֐��D��!��NH��5�����w���or��w��6�$�:�RW��چu5M&�����s��]+��%fr��l��%�i^��3NL��g��\n��K�<�@��[l>�;p�h����6�'H'ā
[��a���mDݠ?��9���2!4�Y����%�,Ikɫߧ3)t~wM)���黣�n;|g;y��%\8m�m��/����	,J?��"U�5㉄tk���y�]�R��[|�	d�k��:��[H��!��g(�`wE5��mݐp����Y�>0W0Z?6{�o�����cxx+�t�ʂ<��]�����=
d�6D�p$�Ёw/�'����VD􊙞���ۚ�?�.؏v����3����Q���q�,�����_ۛA��5�t����3q>�q!IA �`ę�Ȉ�e�v��~~X�uaK�ᨸ�}f6d�V8���Z�A��4I޻��I��.8���L�1��Ǔ,���Л^�,��¥S��JQ�����=� `�U�3V|����#^���]�x��1Vv�2��o�i�y=�w����Y��C;?w��Gaq�pS2��q)=�$E�\LW��JX�j������R����
�
�7�z �2@|8t��5�'�j��}X����sW�ב�(x&�|�O���rFp}�L ��!{\ęu�����	���y#uÖ�HFo���n/<u=�9ӓ�S�tmJ�t���[�8W,��@_��Y0���ы�T��2�4|�#����^G��]8��U��H��J`M-��ʜ�4G���@�����A�X�]`�!iF@-]�lz@�d����ҥ~K4o�.?��׎A岵|��u�3�	�$�I3���D��Ԏ���z'���!���~d ����#I��+�df�L�������i��?~�Do�Z7�� lnr:�'.�0�K.6�p$vuE~p Ek�&?�6r�̘>+�kI��}��>�d����R��A?��byQ��+S��>����$#��_��!��D��� D�>�uΔ��]Z&4]��Ǒ�H[.�9�bz$�΄<\�����6�Zi��6���Y`T9��T��ԖCL�3���L�k�)�`C�Й��O�'ٗ�E�"�-eX? ��?���IhN�5��,:,n^D骬����Hs��8U�99��i��q�[��(CS��V�����lt�W'��/w.���O����`�E荿"�s��J�`͐�����}�k�F#��5�P��	��|�x�\��ϵ�Hp���Wo#��x���u�6�C��wJ�]��W �}��D(���?#��=�	�����û��6���ė0�#�"R9^�� �	���C�<�����xe��m��ST����"�4��Sv��\����ځ�kY%-��@K���C�\(���dxv�?s�����4���fDDn?�$�q�C	������o��`51S"��������������u�����i�_�wT5*�>~�?PK   �^W�e�p  �     jsons/user_defined.json��n�0Ey�J� ;8���&�VQӮ���aKĦ64���{�y4�R�TIw,�=_1w��U�P�Z��[�J.X�l����R���z��f�U��u}�xLF����dɛ|n�k,5o@{�<m�L����`%��6�H�ңyR'��8$���E��aQ��(=L1p�tiܨ�}͓0�+^7�a�s�y~&ޭ�t5#QJ��h	�u���eFC�i�A���I.�`gN+�{�Q1i:�h��<�
*AD]L}�>%� $��p}'�T�><�J3fhc���O��wv�V�xp'׃���zp�a9�>���bx����p��������eǒ+������j�6%̊�R�q��}���ҧK�.��.��'PK   �^Wڮo�  �
            ��    cirkitFile.jsonPK   �^Wġ�e� M� /           ����  images/ff07c967-2774-423d-b98a-e9b309260373.pngPK   �^W�e�p  �             ��N@ jsons/user_defined.jsonPK      �   �A   